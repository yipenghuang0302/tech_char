
module mux ( .data_i({\data_i[31][31] , \data_i[31][30] , \data_i[31][29] , 
        \data_i[31][28] , \data_i[31][27] , \data_i[31][26] , \data_i[31][25] , 
        \data_i[31][24] , \data_i[31][23] , \data_i[31][22] , \data_i[31][21] , 
        \data_i[31][20] , \data_i[31][19] , \data_i[31][18] , \data_i[31][17] , 
        \data_i[31][16] , \data_i[31][15] , \data_i[31][14] , \data_i[31][13] , 
        \data_i[31][12] , \data_i[31][11] , \data_i[31][10] , \data_i[31][9] , 
        \data_i[31][8] , \data_i[31][7] , \data_i[31][6] , \data_i[31][5] , 
        \data_i[31][4] , \data_i[31][3] , \data_i[31][2] , \data_i[31][1] , 
        \data_i[31][0] , \data_i[30][31] , \data_i[30][30] , \data_i[30][29] , 
        \data_i[30][28] , \data_i[30][27] , \data_i[30][26] , \data_i[30][25] , 
        \data_i[30][24] , \data_i[30][23] , \data_i[30][22] , \data_i[30][21] , 
        \data_i[30][20] , \data_i[30][19] , \data_i[30][18] , \data_i[30][17] , 
        \data_i[30][16] , \data_i[30][15] , \data_i[30][14] , \data_i[30][13] , 
        \data_i[30][12] , \data_i[30][11] , \data_i[30][10] , \data_i[30][9] , 
        \data_i[30][8] , \data_i[30][7] , \data_i[30][6] , \data_i[30][5] , 
        \data_i[30][4] , \data_i[30][3] , \data_i[30][2] , \data_i[30][1] , 
        \data_i[30][0] , \data_i[29][31] , \data_i[29][30] , \data_i[29][29] , 
        \data_i[29][28] , \data_i[29][27] , \data_i[29][26] , \data_i[29][25] , 
        \data_i[29][24] , \data_i[29][23] , \data_i[29][22] , \data_i[29][21] , 
        \data_i[29][20] , \data_i[29][19] , \data_i[29][18] , \data_i[29][17] , 
        \data_i[29][16] , \data_i[29][15] , \data_i[29][14] , \data_i[29][13] , 
        \data_i[29][12] , \data_i[29][11] , \data_i[29][10] , \data_i[29][9] , 
        \data_i[29][8] , \data_i[29][7] , \data_i[29][6] , \data_i[29][5] , 
        \data_i[29][4] , \data_i[29][3] , \data_i[29][2] , \data_i[29][1] , 
        \data_i[29][0] , \data_i[28][31] , \data_i[28][30] , \data_i[28][29] , 
        \data_i[28][28] , \data_i[28][27] , \data_i[28][26] , \data_i[28][25] , 
        \data_i[28][24] , \data_i[28][23] , \data_i[28][22] , \data_i[28][21] , 
        \data_i[28][20] , \data_i[28][19] , \data_i[28][18] , \data_i[28][17] , 
        \data_i[28][16] , \data_i[28][15] , \data_i[28][14] , \data_i[28][13] , 
        \data_i[28][12] , \data_i[28][11] , \data_i[28][10] , \data_i[28][9] , 
        \data_i[28][8] , \data_i[28][7] , \data_i[28][6] , \data_i[28][5] , 
        \data_i[28][4] , \data_i[28][3] , \data_i[28][2] , \data_i[28][1] , 
        \data_i[28][0] , \data_i[27][31] , \data_i[27][30] , \data_i[27][29] , 
        \data_i[27][28] , \data_i[27][27] , \data_i[27][26] , \data_i[27][25] , 
        \data_i[27][24] , \data_i[27][23] , \data_i[27][22] , \data_i[27][21] , 
        \data_i[27][20] , \data_i[27][19] , \data_i[27][18] , \data_i[27][17] , 
        \data_i[27][16] , \data_i[27][15] , \data_i[27][14] , \data_i[27][13] , 
        \data_i[27][12] , \data_i[27][11] , \data_i[27][10] , \data_i[27][9] , 
        \data_i[27][8] , \data_i[27][7] , \data_i[27][6] , \data_i[27][5] , 
        \data_i[27][4] , \data_i[27][3] , \data_i[27][2] , \data_i[27][1] , 
        \data_i[27][0] , \data_i[26][31] , \data_i[26][30] , \data_i[26][29] , 
        \data_i[26][28] , \data_i[26][27] , \data_i[26][26] , \data_i[26][25] , 
        \data_i[26][24] , \data_i[26][23] , \data_i[26][22] , \data_i[26][21] , 
        \data_i[26][20] , \data_i[26][19] , \data_i[26][18] , \data_i[26][17] , 
        \data_i[26][16] , \data_i[26][15] , \data_i[26][14] , \data_i[26][13] , 
        \data_i[26][12] , \data_i[26][11] , \data_i[26][10] , \data_i[26][9] , 
        \data_i[26][8] , \data_i[26][7] , \data_i[26][6] , \data_i[26][5] , 
        \data_i[26][4] , \data_i[26][3] , \data_i[26][2] , \data_i[26][1] , 
        \data_i[26][0] , \data_i[25][31] , \data_i[25][30] , \data_i[25][29] , 
        \data_i[25][28] , \data_i[25][27] , \data_i[25][26] , \data_i[25][25] , 
        \data_i[25][24] , \data_i[25][23] , \data_i[25][22] , \data_i[25][21] , 
        \data_i[25][20] , \data_i[25][19] , \data_i[25][18] , \data_i[25][17] , 
        \data_i[25][16] , \data_i[25][15] , \data_i[25][14] , \data_i[25][13] , 
        \data_i[25][12] , \data_i[25][11] , \data_i[25][10] , \data_i[25][9] , 
        \data_i[25][8] , \data_i[25][7] , \data_i[25][6] , \data_i[25][5] , 
        \data_i[25][4] , \data_i[25][3] , \data_i[25][2] , \data_i[25][1] , 
        \data_i[25][0] , \data_i[24][31] , \data_i[24][30] , \data_i[24][29] , 
        \data_i[24][28] , \data_i[24][27] , \data_i[24][26] , \data_i[24][25] , 
        \data_i[24][24] , \data_i[24][23] , \data_i[24][22] , \data_i[24][21] , 
        \data_i[24][20] , \data_i[24][19] , \data_i[24][18] , \data_i[24][17] , 
        \data_i[24][16] , \data_i[24][15] , \data_i[24][14] , \data_i[24][13] , 
        \data_i[24][12] , \data_i[24][11] , \data_i[24][10] , \data_i[24][9] , 
        \data_i[24][8] , \data_i[24][7] , \data_i[24][6] , \data_i[24][5] , 
        \data_i[24][4] , \data_i[24][3] , \data_i[24][2] , \data_i[24][1] , 
        \data_i[24][0] , \data_i[23][31] , \data_i[23][30] , \data_i[23][29] , 
        \data_i[23][28] , \data_i[23][27] , \data_i[23][26] , \data_i[23][25] , 
        \data_i[23][24] , \data_i[23][23] , \data_i[23][22] , \data_i[23][21] , 
        \data_i[23][20] , \data_i[23][19] , \data_i[23][18] , \data_i[23][17] , 
        \data_i[23][16] , \data_i[23][15] , \data_i[23][14] , \data_i[23][13] , 
        \data_i[23][12] , \data_i[23][11] , \data_i[23][10] , \data_i[23][9] , 
        \data_i[23][8] , \data_i[23][7] , \data_i[23][6] , \data_i[23][5] , 
        \data_i[23][4] , \data_i[23][3] , \data_i[23][2] , \data_i[23][1] , 
        \data_i[23][0] , \data_i[22][31] , \data_i[22][30] , \data_i[22][29] , 
        \data_i[22][28] , \data_i[22][27] , \data_i[22][26] , \data_i[22][25] , 
        \data_i[22][24] , \data_i[22][23] , \data_i[22][22] , \data_i[22][21] , 
        \data_i[22][20] , \data_i[22][19] , \data_i[22][18] , \data_i[22][17] , 
        \data_i[22][16] , \data_i[22][15] , \data_i[22][14] , \data_i[22][13] , 
        \data_i[22][12] , \data_i[22][11] , \data_i[22][10] , \data_i[22][9] , 
        \data_i[22][8] , \data_i[22][7] , \data_i[22][6] , \data_i[22][5] , 
        \data_i[22][4] , \data_i[22][3] , \data_i[22][2] , \data_i[22][1] , 
        \data_i[22][0] , \data_i[21][31] , \data_i[21][30] , \data_i[21][29] , 
        \data_i[21][28] , \data_i[21][27] , \data_i[21][26] , \data_i[21][25] , 
        \data_i[21][24] , \data_i[21][23] , \data_i[21][22] , \data_i[21][21] , 
        \data_i[21][20] , \data_i[21][19] , \data_i[21][18] , \data_i[21][17] , 
        \data_i[21][16] , \data_i[21][15] , \data_i[21][14] , \data_i[21][13] , 
        \data_i[21][12] , \data_i[21][11] , \data_i[21][10] , \data_i[21][9] , 
        \data_i[21][8] , \data_i[21][7] , \data_i[21][6] , \data_i[21][5] , 
        \data_i[21][4] , \data_i[21][3] , \data_i[21][2] , \data_i[21][1] , 
        \data_i[21][0] , \data_i[20][31] , \data_i[20][30] , \data_i[20][29] , 
        \data_i[20][28] , \data_i[20][27] , \data_i[20][26] , \data_i[20][25] , 
        \data_i[20][24] , \data_i[20][23] , \data_i[20][22] , \data_i[20][21] , 
        \data_i[20][20] , \data_i[20][19] , \data_i[20][18] , \data_i[20][17] , 
        \data_i[20][16] , \data_i[20][15] , \data_i[20][14] , \data_i[20][13] , 
        \data_i[20][12] , \data_i[20][11] , \data_i[20][10] , \data_i[20][9] , 
        \data_i[20][8] , \data_i[20][7] , \data_i[20][6] , \data_i[20][5] , 
        \data_i[20][4] , \data_i[20][3] , \data_i[20][2] , \data_i[20][1] , 
        \data_i[20][0] , \data_i[19][31] , \data_i[19][30] , \data_i[19][29] , 
        \data_i[19][28] , \data_i[19][27] , \data_i[19][26] , \data_i[19][25] , 
        \data_i[19][24] , \data_i[19][23] , \data_i[19][22] , \data_i[19][21] , 
        \data_i[19][20] , \data_i[19][19] , \data_i[19][18] , \data_i[19][17] , 
        \data_i[19][16] , \data_i[19][15] , \data_i[19][14] , \data_i[19][13] , 
        \data_i[19][12] , \data_i[19][11] , \data_i[19][10] , \data_i[19][9] , 
        \data_i[19][8] , \data_i[19][7] , \data_i[19][6] , \data_i[19][5] , 
        \data_i[19][4] , \data_i[19][3] , \data_i[19][2] , \data_i[19][1] , 
        \data_i[19][0] , \data_i[18][31] , \data_i[18][30] , \data_i[18][29] , 
        \data_i[18][28] , \data_i[18][27] , \data_i[18][26] , \data_i[18][25] , 
        \data_i[18][24] , \data_i[18][23] , \data_i[18][22] , \data_i[18][21] , 
        \data_i[18][20] , \data_i[18][19] , \data_i[18][18] , \data_i[18][17] , 
        \data_i[18][16] , \data_i[18][15] , \data_i[18][14] , \data_i[18][13] , 
        \data_i[18][12] , \data_i[18][11] , \data_i[18][10] , \data_i[18][9] , 
        \data_i[18][8] , \data_i[18][7] , \data_i[18][6] , \data_i[18][5] , 
        \data_i[18][4] , \data_i[18][3] , \data_i[18][2] , \data_i[18][1] , 
        \data_i[18][0] , \data_i[17][31] , \data_i[17][30] , \data_i[17][29] , 
        \data_i[17][28] , \data_i[17][27] , \data_i[17][26] , \data_i[17][25] , 
        \data_i[17][24] , \data_i[17][23] , \data_i[17][22] , \data_i[17][21] , 
        \data_i[17][20] , \data_i[17][19] , \data_i[17][18] , \data_i[17][17] , 
        \data_i[17][16] , \data_i[17][15] , \data_i[17][14] , \data_i[17][13] , 
        \data_i[17][12] , \data_i[17][11] , \data_i[17][10] , \data_i[17][9] , 
        \data_i[17][8] , \data_i[17][7] , \data_i[17][6] , \data_i[17][5] , 
        \data_i[17][4] , \data_i[17][3] , \data_i[17][2] , \data_i[17][1] , 
        \data_i[17][0] , \data_i[16][31] , \data_i[16][30] , \data_i[16][29] , 
        \data_i[16][28] , \data_i[16][27] , \data_i[16][26] , \data_i[16][25] , 
        \data_i[16][24] , \data_i[16][23] , \data_i[16][22] , \data_i[16][21] , 
        \data_i[16][20] , \data_i[16][19] , \data_i[16][18] , \data_i[16][17] , 
        \data_i[16][16] , \data_i[16][15] , \data_i[16][14] , \data_i[16][13] , 
        \data_i[16][12] , \data_i[16][11] , \data_i[16][10] , \data_i[16][9] , 
        \data_i[16][8] , \data_i[16][7] , \data_i[16][6] , \data_i[16][5] , 
        \data_i[16][4] , \data_i[16][3] , \data_i[16][2] , \data_i[16][1] , 
        \data_i[16][0] , \data_i[15][31] , \data_i[15][30] , \data_i[15][29] , 
        \data_i[15][28] , \data_i[15][27] , \data_i[15][26] , \data_i[15][25] , 
        \data_i[15][24] , \data_i[15][23] , \data_i[15][22] , \data_i[15][21] , 
        \data_i[15][20] , \data_i[15][19] , \data_i[15][18] , \data_i[15][17] , 
        \data_i[15][16] , \data_i[15][15] , \data_i[15][14] , \data_i[15][13] , 
        \data_i[15][12] , \data_i[15][11] , \data_i[15][10] , \data_i[15][9] , 
        \data_i[15][8] , \data_i[15][7] , \data_i[15][6] , \data_i[15][5] , 
        \data_i[15][4] , \data_i[15][3] , \data_i[15][2] , \data_i[15][1] , 
        \data_i[15][0] , \data_i[14][31] , \data_i[14][30] , \data_i[14][29] , 
        \data_i[14][28] , \data_i[14][27] , \data_i[14][26] , \data_i[14][25] , 
        \data_i[14][24] , \data_i[14][23] , \data_i[14][22] , \data_i[14][21] , 
        \data_i[14][20] , \data_i[14][19] , \data_i[14][18] , \data_i[14][17] , 
        \data_i[14][16] , \data_i[14][15] , \data_i[14][14] , \data_i[14][13] , 
        \data_i[14][12] , \data_i[14][11] , \data_i[14][10] , \data_i[14][9] , 
        \data_i[14][8] , \data_i[14][7] , \data_i[14][6] , \data_i[14][5] , 
        \data_i[14][4] , \data_i[14][3] , \data_i[14][2] , \data_i[14][1] , 
        \data_i[14][0] , \data_i[13][31] , \data_i[13][30] , \data_i[13][29] , 
        \data_i[13][28] , \data_i[13][27] , \data_i[13][26] , \data_i[13][25] , 
        \data_i[13][24] , \data_i[13][23] , \data_i[13][22] , \data_i[13][21] , 
        \data_i[13][20] , \data_i[13][19] , \data_i[13][18] , \data_i[13][17] , 
        \data_i[13][16] , \data_i[13][15] , \data_i[13][14] , \data_i[13][13] , 
        \data_i[13][12] , \data_i[13][11] , \data_i[13][10] , \data_i[13][9] , 
        \data_i[13][8] , \data_i[13][7] , \data_i[13][6] , \data_i[13][5] , 
        \data_i[13][4] , \data_i[13][3] , \data_i[13][2] , \data_i[13][1] , 
        \data_i[13][0] , \data_i[12][31] , \data_i[12][30] , \data_i[12][29] , 
        \data_i[12][28] , \data_i[12][27] , \data_i[12][26] , \data_i[12][25] , 
        \data_i[12][24] , \data_i[12][23] , \data_i[12][22] , \data_i[12][21] , 
        \data_i[12][20] , \data_i[12][19] , \data_i[12][18] , \data_i[12][17] , 
        \data_i[12][16] , \data_i[12][15] , \data_i[12][14] , \data_i[12][13] , 
        \data_i[12][12] , \data_i[12][11] , \data_i[12][10] , \data_i[12][9] , 
        \data_i[12][8] , \data_i[12][7] , \data_i[12][6] , \data_i[12][5] , 
        \data_i[12][4] , \data_i[12][3] , \data_i[12][2] , \data_i[12][1] , 
        \data_i[12][0] , \data_i[11][31] , \data_i[11][30] , \data_i[11][29] , 
        \data_i[11][28] , \data_i[11][27] , \data_i[11][26] , \data_i[11][25] , 
        \data_i[11][24] , \data_i[11][23] , \data_i[11][22] , \data_i[11][21] , 
        \data_i[11][20] , \data_i[11][19] , \data_i[11][18] , \data_i[11][17] , 
        \data_i[11][16] , \data_i[11][15] , \data_i[11][14] , \data_i[11][13] , 
        \data_i[11][12] , \data_i[11][11] , \data_i[11][10] , \data_i[11][9] , 
        \data_i[11][8] , \data_i[11][7] , \data_i[11][6] , \data_i[11][5] , 
        \data_i[11][4] , \data_i[11][3] , \data_i[11][2] , \data_i[11][1] , 
        \data_i[11][0] , \data_i[10][31] , \data_i[10][30] , \data_i[10][29] , 
        \data_i[10][28] , \data_i[10][27] , \data_i[10][26] , \data_i[10][25] , 
        \data_i[10][24] , \data_i[10][23] , \data_i[10][22] , \data_i[10][21] , 
        \data_i[10][20] , \data_i[10][19] , \data_i[10][18] , \data_i[10][17] , 
        \data_i[10][16] , \data_i[10][15] , \data_i[10][14] , \data_i[10][13] , 
        \data_i[10][12] , \data_i[10][11] , \data_i[10][10] , \data_i[10][9] , 
        \data_i[10][8] , \data_i[10][7] , \data_i[10][6] , \data_i[10][5] , 
        \data_i[10][4] , \data_i[10][3] , \data_i[10][2] , \data_i[10][1] , 
        \data_i[10][0] , \data_i[9][31] , \data_i[9][30] , \data_i[9][29] , 
        \data_i[9][28] , \data_i[9][27] , \data_i[9][26] , \data_i[9][25] , 
        \data_i[9][24] , \data_i[9][23] , \data_i[9][22] , \data_i[9][21] , 
        \data_i[9][20] , \data_i[9][19] , \data_i[9][18] , \data_i[9][17] , 
        \data_i[9][16] , \data_i[9][15] , \data_i[9][14] , \data_i[9][13] , 
        \data_i[9][12] , \data_i[9][11] , \data_i[9][10] , \data_i[9][9] , 
        \data_i[9][8] , \data_i[9][7] , \data_i[9][6] , \data_i[9][5] , 
        \data_i[9][4] , \data_i[9][3] , \data_i[9][2] , \data_i[9][1] , 
        \data_i[9][0] , \data_i[8][31] , \data_i[8][30] , \data_i[8][29] , 
        \data_i[8][28] , \data_i[8][27] , \data_i[8][26] , \data_i[8][25] , 
        \data_i[8][24] , \data_i[8][23] , \data_i[8][22] , \data_i[8][21] , 
        \data_i[8][20] , \data_i[8][19] , \data_i[8][18] , \data_i[8][17] , 
        \data_i[8][16] , \data_i[8][15] , \data_i[8][14] , \data_i[8][13] , 
        \data_i[8][12] , \data_i[8][11] , \data_i[8][10] , \data_i[8][9] , 
        \data_i[8][8] , \data_i[8][7] , \data_i[8][6] , \data_i[8][5] , 
        \data_i[8][4] , \data_i[8][3] , \data_i[8][2] , \data_i[8][1] , 
        \data_i[8][0] , \data_i[7][31] , \data_i[7][30] , \data_i[7][29] , 
        \data_i[7][28] , \data_i[7][27] , \data_i[7][26] , \data_i[7][25] , 
        \data_i[7][24] , \data_i[7][23] , \data_i[7][22] , \data_i[7][21] , 
        \data_i[7][20] , \data_i[7][19] , \data_i[7][18] , \data_i[7][17] , 
        \data_i[7][16] , \data_i[7][15] , \data_i[7][14] , \data_i[7][13] , 
        \data_i[7][12] , \data_i[7][11] , \data_i[7][10] , \data_i[7][9] , 
        \data_i[7][8] , \data_i[7][7] , \data_i[7][6] , \data_i[7][5] , 
        \data_i[7][4] , \data_i[7][3] , \data_i[7][2] , \data_i[7][1] , 
        \data_i[7][0] , \data_i[6][31] , \data_i[6][30] , \data_i[6][29] , 
        \data_i[6][28] , \data_i[6][27] , \data_i[6][26] , \data_i[6][25] , 
        \data_i[6][24] , \data_i[6][23] , \data_i[6][22] , \data_i[6][21] , 
        \data_i[6][20] , \data_i[6][19] , \data_i[6][18] , \data_i[6][17] , 
        \data_i[6][16] , \data_i[6][15] , \data_i[6][14] , \data_i[6][13] , 
        \data_i[6][12] , \data_i[6][11] , \data_i[6][10] , \data_i[6][9] , 
        \data_i[6][8] , \data_i[6][7] , \data_i[6][6] , \data_i[6][5] , 
        \data_i[6][4] , \data_i[6][3] , \data_i[6][2] , \data_i[6][1] , 
        \data_i[6][0] , \data_i[5][31] , \data_i[5][30] , \data_i[5][29] , 
        \data_i[5][28] , \data_i[5][27] , \data_i[5][26] , \data_i[5][25] , 
        \data_i[5][24] , \data_i[5][23] , \data_i[5][22] , \data_i[5][21] , 
        \data_i[5][20] , \data_i[5][19] , \data_i[5][18] , \data_i[5][17] , 
        \data_i[5][16] , \data_i[5][15] , \data_i[5][14] , \data_i[5][13] , 
        \data_i[5][12] , \data_i[5][11] , \data_i[5][10] , \data_i[5][9] , 
        \data_i[5][8] , \data_i[5][7] , \data_i[5][6] , \data_i[5][5] , 
        \data_i[5][4] , \data_i[5][3] , \data_i[5][2] , \data_i[5][1] , 
        \data_i[5][0] , \data_i[4][31] , \data_i[4][30] , \data_i[4][29] , 
        \data_i[4][28] , \data_i[4][27] , \data_i[4][26] , \data_i[4][25] , 
        \data_i[4][24] , \data_i[4][23] , \data_i[4][22] , \data_i[4][21] , 
        \data_i[4][20] , \data_i[4][19] , \data_i[4][18] , \data_i[4][17] , 
        \data_i[4][16] , \data_i[4][15] , \data_i[4][14] , \data_i[4][13] , 
        \data_i[4][12] , \data_i[4][11] , \data_i[4][10] , \data_i[4][9] , 
        \data_i[4][8] , \data_i[4][7] , \data_i[4][6] , \data_i[4][5] , 
        \data_i[4][4] , \data_i[4][3] , \data_i[4][2] , \data_i[4][1] , 
        \data_i[4][0] , \data_i[3][31] , \data_i[3][30] , \data_i[3][29] , 
        \data_i[3][28] , \data_i[3][27] , \data_i[3][26] , \data_i[3][25] , 
        \data_i[3][24] , \data_i[3][23] , \data_i[3][22] , \data_i[3][21] , 
        \data_i[3][20] , \data_i[3][19] , \data_i[3][18] , \data_i[3][17] , 
        \data_i[3][16] , \data_i[3][15] , \data_i[3][14] , \data_i[3][13] , 
        \data_i[3][12] , \data_i[3][11] , \data_i[3][10] , \data_i[3][9] , 
        \data_i[3][8] , \data_i[3][7] , \data_i[3][6] , \data_i[3][5] , 
        \data_i[3][4] , \data_i[3][3] , \data_i[3][2] , \data_i[3][1] , 
        \data_i[3][0] , \data_i[2][31] , \data_i[2][30] , \data_i[2][29] , 
        \data_i[2][28] , \data_i[2][27] , \data_i[2][26] , \data_i[2][25] , 
        \data_i[2][24] , \data_i[2][23] , \data_i[2][22] , \data_i[2][21] , 
        \data_i[2][20] , \data_i[2][19] , \data_i[2][18] , \data_i[2][17] , 
        \data_i[2][16] , \data_i[2][15] , \data_i[2][14] , \data_i[2][13] , 
        \data_i[2][12] , \data_i[2][11] , \data_i[2][10] , \data_i[2][9] , 
        \data_i[2][8] , \data_i[2][7] , \data_i[2][6] , \data_i[2][5] , 
        \data_i[2][4] , \data_i[2][3] , \data_i[2][2] , \data_i[2][1] , 
        \data_i[2][0] , \data_i[1][31] , \data_i[1][30] , \data_i[1][29] , 
        \data_i[1][28] , \data_i[1][27] , \data_i[1][26] , \data_i[1][25] , 
        \data_i[1][24] , \data_i[1][23] , \data_i[1][22] , \data_i[1][21] , 
        \data_i[1][20] , \data_i[1][19] , \data_i[1][18] , \data_i[1][17] , 
        \data_i[1][16] , \data_i[1][15] , \data_i[1][14] , \data_i[1][13] , 
        \data_i[1][12] , \data_i[1][11] , \data_i[1][10] , \data_i[1][9] , 
        \data_i[1][8] , \data_i[1][7] , \data_i[1][6] , \data_i[1][5] , 
        \data_i[1][4] , \data_i[1][3] , \data_i[1][2] , \data_i[1][1] , 
        \data_i[1][0] , \data_i[0][31] , \data_i[0][30] , \data_i[0][29] , 
        \data_i[0][28] , \data_i[0][27] , \data_i[0][26] , \data_i[0][25] , 
        \data_i[0][24] , \data_i[0][23] , \data_i[0][22] , \data_i[0][21] , 
        \data_i[0][20] , \data_i[0][19] , \data_i[0][18] , \data_i[0][17] , 
        \data_i[0][16] , \data_i[0][15] , \data_i[0][14] , \data_i[0][13] , 
        \data_i[0][12] , \data_i[0][11] , \data_i[0][10] , \data_i[0][9] , 
        \data_i[0][8] , \data_i[0][7] , \data_i[0][6] , \data_i[0][5] , 
        \data_i[0][4] , \data_i[0][3] , \data_i[0][2] , \data_i[0][1] , 
        \data_i[0][0] }), select_i, data_o );
  input [4:0] select_i;
  output [31:0] data_o;
  input \data_i[31][31] , \data_i[31][30] , \data_i[31][29] , \data_i[31][28] ,
         \data_i[31][27] , \data_i[31][26] , \data_i[31][25] ,
         \data_i[31][24] , \data_i[31][23] , \data_i[31][22] ,
         \data_i[31][21] , \data_i[31][20] , \data_i[31][19] ,
         \data_i[31][18] , \data_i[31][17] , \data_i[31][16] ,
         \data_i[31][15] , \data_i[31][14] , \data_i[31][13] ,
         \data_i[31][12] , \data_i[31][11] , \data_i[31][10] , \data_i[31][9] ,
         \data_i[31][8] , \data_i[31][7] , \data_i[31][6] , \data_i[31][5] ,
         \data_i[31][4] , \data_i[31][3] , \data_i[31][2] , \data_i[31][1] ,
         \data_i[31][0] , \data_i[30][31] , \data_i[30][30] , \data_i[30][29] ,
         \data_i[30][28] , \data_i[30][27] , \data_i[30][26] ,
         \data_i[30][25] , \data_i[30][24] , \data_i[30][23] ,
         \data_i[30][22] , \data_i[30][21] , \data_i[30][20] ,
         \data_i[30][19] , \data_i[30][18] , \data_i[30][17] ,
         \data_i[30][16] , \data_i[30][15] , \data_i[30][14] ,
         \data_i[30][13] , \data_i[30][12] , \data_i[30][11] ,
         \data_i[30][10] , \data_i[30][9] , \data_i[30][8] , \data_i[30][7] ,
         \data_i[30][6] , \data_i[30][5] , \data_i[30][4] , \data_i[30][3] ,
         \data_i[30][2] , \data_i[30][1] , \data_i[30][0] , \data_i[29][31] ,
         \data_i[29][30] , \data_i[29][29] , \data_i[29][28] ,
         \data_i[29][27] , \data_i[29][26] , \data_i[29][25] ,
         \data_i[29][24] , \data_i[29][23] , \data_i[29][22] ,
         \data_i[29][21] , \data_i[29][20] , \data_i[29][19] ,
         \data_i[29][18] , \data_i[29][17] , \data_i[29][16] ,
         \data_i[29][15] , \data_i[29][14] , \data_i[29][13] ,
         \data_i[29][12] , \data_i[29][11] , \data_i[29][10] , \data_i[29][9] ,
         \data_i[29][8] , \data_i[29][7] , \data_i[29][6] , \data_i[29][5] ,
         \data_i[29][4] , \data_i[29][3] , \data_i[29][2] , \data_i[29][1] ,
         \data_i[29][0] , \data_i[28][31] , \data_i[28][30] , \data_i[28][29] ,
         \data_i[28][28] , \data_i[28][27] , \data_i[28][26] ,
         \data_i[28][25] , \data_i[28][24] , \data_i[28][23] ,
         \data_i[28][22] , \data_i[28][21] , \data_i[28][20] ,
         \data_i[28][19] , \data_i[28][18] , \data_i[28][17] ,
         \data_i[28][16] , \data_i[28][15] , \data_i[28][14] ,
         \data_i[28][13] , \data_i[28][12] , \data_i[28][11] ,
         \data_i[28][10] , \data_i[28][9] , \data_i[28][8] , \data_i[28][7] ,
         \data_i[28][6] , \data_i[28][5] , \data_i[28][4] , \data_i[28][3] ,
         \data_i[28][2] , \data_i[28][1] , \data_i[28][0] , \data_i[27][31] ,
         \data_i[27][30] , \data_i[27][29] , \data_i[27][28] ,
         \data_i[27][27] , \data_i[27][26] , \data_i[27][25] ,
         \data_i[27][24] , \data_i[27][23] , \data_i[27][22] ,
         \data_i[27][21] , \data_i[27][20] , \data_i[27][19] ,
         \data_i[27][18] , \data_i[27][17] , \data_i[27][16] ,
         \data_i[27][15] , \data_i[27][14] , \data_i[27][13] ,
         \data_i[27][12] , \data_i[27][11] , \data_i[27][10] , \data_i[27][9] ,
         \data_i[27][8] , \data_i[27][7] , \data_i[27][6] , \data_i[27][5] ,
         \data_i[27][4] , \data_i[27][3] , \data_i[27][2] , \data_i[27][1] ,
         \data_i[27][0] , \data_i[26][31] , \data_i[26][30] , \data_i[26][29] ,
         \data_i[26][28] , \data_i[26][27] , \data_i[26][26] ,
         \data_i[26][25] , \data_i[26][24] , \data_i[26][23] ,
         \data_i[26][22] , \data_i[26][21] , \data_i[26][20] ,
         \data_i[26][19] , \data_i[26][18] , \data_i[26][17] ,
         \data_i[26][16] , \data_i[26][15] , \data_i[26][14] ,
         \data_i[26][13] , \data_i[26][12] , \data_i[26][11] ,
         \data_i[26][10] , \data_i[26][9] , \data_i[26][8] , \data_i[26][7] ,
         \data_i[26][6] , \data_i[26][5] , \data_i[26][4] , \data_i[26][3] ,
         \data_i[26][2] , \data_i[26][1] , \data_i[26][0] , \data_i[25][31] ,
         \data_i[25][30] , \data_i[25][29] , \data_i[25][28] ,
         \data_i[25][27] , \data_i[25][26] , \data_i[25][25] ,
         \data_i[25][24] , \data_i[25][23] , \data_i[25][22] ,
         \data_i[25][21] , \data_i[25][20] , \data_i[25][19] ,
         \data_i[25][18] , \data_i[25][17] , \data_i[25][16] ,
         \data_i[25][15] , \data_i[25][14] , \data_i[25][13] ,
         \data_i[25][12] , \data_i[25][11] , \data_i[25][10] , \data_i[25][9] ,
         \data_i[25][8] , \data_i[25][7] , \data_i[25][6] , \data_i[25][5] ,
         \data_i[25][4] , \data_i[25][3] , \data_i[25][2] , \data_i[25][1] ,
         \data_i[25][0] , \data_i[24][31] , \data_i[24][30] , \data_i[24][29] ,
         \data_i[24][28] , \data_i[24][27] , \data_i[24][26] ,
         \data_i[24][25] , \data_i[24][24] , \data_i[24][23] ,
         \data_i[24][22] , \data_i[24][21] , \data_i[24][20] ,
         \data_i[24][19] , \data_i[24][18] , \data_i[24][17] ,
         \data_i[24][16] , \data_i[24][15] , \data_i[24][14] ,
         \data_i[24][13] , \data_i[24][12] , \data_i[24][11] ,
         \data_i[24][10] , \data_i[24][9] , \data_i[24][8] , \data_i[24][7] ,
         \data_i[24][6] , \data_i[24][5] , \data_i[24][4] , \data_i[24][3] ,
         \data_i[24][2] , \data_i[24][1] , \data_i[24][0] , \data_i[23][31] ,
         \data_i[23][30] , \data_i[23][29] , \data_i[23][28] ,
         \data_i[23][27] , \data_i[23][26] , \data_i[23][25] ,
         \data_i[23][24] , \data_i[23][23] , \data_i[23][22] ,
         \data_i[23][21] , \data_i[23][20] , \data_i[23][19] ,
         \data_i[23][18] , \data_i[23][17] , \data_i[23][16] ,
         \data_i[23][15] , \data_i[23][14] , \data_i[23][13] ,
         \data_i[23][12] , \data_i[23][11] , \data_i[23][10] , \data_i[23][9] ,
         \data_i[23][8] , \data_i[23][7] , \data_i[23][6] , \data_i[23][5] ,
         \data_i[23][4] , \data_i[23][3] , \data_i[23][2] , \data_i[23][1] ,
         \data_i[23][0] , \data_i[22][31] , \data_i[22][30] , \data_i[22][29] ,
         \data_i[22][28] , \data_i[22][27] , \data_i[22][26] ,
         \data_i[22][25] , \data_i[22][24] , \data_i[22][23] ,
         \data_i[22][22] , \data_i[22][21] , \data_i[22][20] ,
         \data_i[22][19] , \data_i[22][18] , \data_i[22][17] ,
         \data_i[22][16] , \data_i[22][15] , \data_i[22][14] ,
         \data_i[22][13] , \data_i[22][12] , \data_i[22][11] ,
         \data_i[22][10] , \data_i[22][9] , \data_i[22][8] , \data_i[22][7] ,
         \data_i[22][6] , \data_i[22][5] , \data_i[22][4] , \data_i[22][3] ,
         \data_i[22][2] , \data_i[22][1] , \data_i[22][0] , \data_i[21][31] ,
         \data_i[21][30] , \data_i[21][29] , \data_i[21][28] ,
         \data_i[21][27] , \data_i[21][26] , \data_i[21][25] ,
         \data_i[21][24] , \data_i[21][23] , \data_i[21][22] ,
         \data_i[21][21] , \data_i[21][20] , \data_i[21][19] ,
         \data_i[21][18] , \data_i[21][17] , \data_i[21][16] ,
         \data_i[21][15] , \data_i[21][14] , \data_i[21][13] ,
         \data_i[21][12] , \data_i[21][11] , \data_i[21][10] , \data_i[21][9] ,
         \data_i[21][8] , \data_i[21][7] , \data_i[21][6] , \data_i[21][5] ,
         \data_i[21][4] , \data_i[21][3] , \data_i[21][2] , \data_i[21][1] ,
         \data_i[21][0] , \data_i[20][31] , \data_i[20][30] , \data_i[20][29] ,
         \data_i[20][28] , \data_i[20][27] , \data_i[20][26] ,
         \data_i[20][25] , \data_i[20][24] , \data_i[20][23] ,
         \data_i[20][22] , \data_i[20][21] , \data_i[20][20] ,
         \data_i[20][19] , \data_i[20][18] , \data_i[20][17] ,
         \data_i[20][16] , \data_i[20][15] , \data_i[20][14] ,
         \data_i[20][13] , \data_i[20][12] , \data_i[20][11] ,
         \data_i[20][10] , \data_i[20][9] , \data_i[20][8] , \data_i[20][7] ,
         \data_i[20][6] , \data_i[20][5] , \data_i[20][4] , \data_i[20][3] ,
         \data_i[20][2] , \data_i[20][1] , \data_i[20][0] , \data_i[19][31] ,
         \data_i[19][30] , \data_i[19][29] , \data_i[19][28] ,
         \data_i[19][27] , \data_i[19][26] , \data_i[19][25] ,
         \data_i[19][24] , \data_i[19][23] , \data_i[19][22] ,
         \data_i[19][21] , \data_i[19][20] , \data_i[19][19] ,
         \data_i[19][18] , \data_i[19][17] , \data_i[19][16] ,
         \data_i[19][15] , \data_i[19][14] , \data_i[19][13] ,
         \data_i[19][12] , \data_i[19][11] , \data_i[19][10] , \data_i[19][9] ,
         \data_i[19][8] , \data_i[19][7] , \data_i[19][6] , \data_i[19][5] ,
         \data_i[19][4] , \data_i[19][3] , \data_i[19][2] , \data_i[19][1] ,
         \data_i[19][0] , \data_i[18][31] , \data_i[18][30] , \data_i[18][29] ,
         \data_i[18][28] , \data_i[18][27] , \data_i[18][26] ,
         \data_i[18][25] , \data_i[18][24] , \data_i[18][23] ,
         \data_i[18][22] , \data_i[18][21] , \data_i[18][20] ,
         \data_i[18][19] , \data_i[18][18] , \data_i[18][17] ,
         \data_i[18][16] , \data_i[18][15] , \data_i[18][14] ,
         \data_i[18][13] , \data_i[18][12] , \data_i[18][11] ,
         \data_i[18][10] , \data_i[18][9] , \data_i[18][8] , \data_i[18][7] ,
         \data_i[18][6] , \data_i[18][5] , \data_i[18][4] , \data_i[18][3] ,
         \data_i[18][2] , \data_i[18][1] , \data_i[18][0] , \data_i[17][31] ,
         \data_i[17][30] , \data_i[17][29] , \data_i[17][28] ,
         \data_i[17][27] , \data_i[17][26] , \data_i[17][25] ,
         \data_i[17][24] , \data_i[17][23] , \data_i[17][22] ,
         \data_i[17][21] , \data_i[17][20] , \data_i[17][19] ,
         \data_i[17][18] , \data_i[17][17] , \data_i[17][16] ,
         \data_i[17][15] , \data_i[17][14] , \data_i[17][13] ,
         \data_i[17][12] , \data_i[17][11] , \data_i[17][10] , \data_i[17][9] ,
         \data_i[17][8] , \data_i[17][7] , \data_i[17][6] , \data_i[17][5] ,
         \data_i[17][4] , \data_i[17][3] , \data_i[17][2] , \data_i[17][1] ,
         \data_i[17][0] , \data_i[16][31] , \data_i[16][30] , \data_i[16][29] ,
         \data_i[16][28] , \data_i[16][27] , \data_i[16][26] ,
         \data_i[16][25] , \data_i[16][24] , \data_i[16][23] ,
         \data_i[16][22] , \data_i[16][21] , \data_i[16][20] ,
         \data_i[16][19] , \data_i[16][18] , \data_i[16][17] ,
         \data_i[16][16] , \data_i[16][15] , \data_i[16][14] ,
         \data_i[16][13] , \data_i[16][12] , \data_i[16][11] ,
         \data_i[16][10] , \data_i[16][9] , \data_i[16][8] , \data_i[16][7] ,
         \data_i[16][6] , \data_i[16][5] , \data_i[16][4] , \data_i[16][3] ,
         \data_i[16][2] , \data_i[16][1] , \data_i[16][0] , \data_i[15][31] ,
         \data_i[15][30] , \data_i[15][29] , \data_i[15][28] ,
         \data_i[15][27] , \data_i[15][26] , \data_i[15][25] ,
         \data_i[15][24] , \data_i[15][23] , \data_i[15][22] ,
         \data_i[15][21] , \data_i[15][20] , \data_i[15][19] ,
         \data_i[15][18] , \data_i[15][17] , \data_i[15][16] ,
         \data_i[15][15] , \data_i[15][14] , \data_i[15][13] ,
         \data_i[15][12] , \data_i[15][11] , \data_i[15][10] , \data_i[15][9] ,
         \data_i[15][8] , \data_i[15][7] , \data_i[15][6] , \data_i[15][5] ,
         \data_i[15][4] , \data_i[15][3] , \data_i[15][2] , \data_i[15][1] ,
         \data_i[15][0] , \data_i[14][31] , \data_i[14][30] , \data_i[14][29] ,
         \data_i[14][28] , \data_i[14][27] , \data_i[14][26] ,
         \data_i[14][25] , \data_i[14][24] , \data_i[14][23] ,
         \data_i[14][22] , \data_i[14][21] , \data_i[14][20] ,
         \data_i[14][19] , \data_i[14][18] , \data_i[14][17] ,
         \data_i[14][16] , \data_i[14][15] , \data_i[14][14] ,
         \data_i[14][13] , \data_i[14][12] , \data_i[14][11] ,
         \data_i[14][10] , \data_i[14][9] , \data_i[14][8] , \data_i[14][7] ,
         \data_i[14][6] , \data_i[14][5] , \data_i[14][4] , \data_i[14][3] ,
         \data_i[14][2] , \data_i[14][1] , \data_i[14][0] , \data_i[13][31] ,
         \data_i[13][30] , \data_i[13][29] , \data_i[13][28] ,
         \data_i[13][27] , \data_i[13][26] , \data_i[13][25] ,
         \data_i[13][24] , \data_i[13][23] , \data_i[13][22] ,
         \data_i[13][21] , \data_i[13][20] , \data_i[13][19] ,
         \data_i[13][18] , \data_i[13][17] , \data_i[13][16] ,
         \data_i[13][15] , \data_i[13][14] , \data_i[13][13] ,
         \data_i[13][12] , \data_i[13][11] , \data_i[13][10] , \data_i[13][9] ,
         \data_i[13][8] , \data_i[13][7] , \data_i[13][6] , \data_i[13][5] ,
         \data_i[13][4] , \data_i[13][3] , \data_i[13][2] , \data_i[13][1] ,
         \data_i[13][0] , \data_i[12][31] , \data_i[12][30] , \data_i[12][29] ,
         \data_i[12][28] , \data_i[12][27] , \data_i[12][26] ,
         \data_i[12][25] , \data_i[12][24] , \data_i[12][23] ,
         \data_i[12][22] , \data_i[12][21] , \data_i[12][20] ,
         \data_i[12][19] , \data_i[12][18] , \data_i[12][17] ,
         \data_i[12][16] , \data_i[12][15] , \data_i[12][14] ,
         \data_i[12][13] , \data_i[12][12] , \data_i[12][11] ,
         \data_i[12][10] , \data_i[12][9] , \data_i[12][8] , \data_i[12][7] ,
         \data_i[12][6] , \data_i[12][5] , \data_i[12][4] , \data_i[12][3] ,
         \data_i[12][2] , \data_i[12][1] , \data_i[12][0] , \data_i[11][31] ,
         \data_i[11][30] , \data_i[11][29] , \data_i[11][28] ,
         \data_i[11][27] , \data_i[11][26] , \data_i[11][25] ,
         \data_i[11][24] , \data_i[11][23] , \data_i[11][22] ,
         \data_i[11][21] , \data_i[11][20] , \data_i[11][19] ,
         \data_i[11][18] , \data_i[11][17] , \data_i[11][16] ,
         \data_i[11][15] , \data_i[11][14] , \data_i[11][13] ,
         \data_i[11][12] , \data_i[11][11] , \data_i[11][10] , \data_i[11][9] ,
         \data_i[11][8] , \data_i[11][7] , \data_i[11][6] , \data_i[11][5] ,
         \data_i[11][4] , \data_i[11][3] , \data_i[11][2] , \data_i[11][1] ,
         \data_i[11][0] , \data_i[10][31] , \data_i[10][30] , \data_i[10][29] ,
         \data_i[10][28] , \data_i[10][27] , \data_i[10][26] ,
         \data_i[10][25] , \data_i[10][24] , \data_i[10][23] ,
         \data_i[10][22] , \data_i[10][21] , \data_i[10][20] ,
         \data_i[10][19] , \data_i[10][18] , \data_i[10][17] ,
         \data_i[10][16] , \data_i[10][15] , \data_i[10][14] ,
         \data_i[10][13] , \data_i[10][12] , \data_i[10][11] ,
         \data_i[10][10] , \data_i[10][9] , \data_i[10][8] , \data_i[10][7] ,
         \data_i[10][6] , \data_i[10][5] , \data_i[10][4] , \data_i[10][3] ,
         \data_i[10][2] , \data_i[10][1] , \data_i[10][0] , \data_i[9][31] ,
         \data_i[9][30] , \data_i[9][29] , \data_i[9][28] , \data_i[9][27] ,
         \data_i[9][26] , \data_i[9][25] , \data_i[9][24] , \data_i[9][23] ,
         \data_i[9][22] , \data_i[9][21] , \data_i[9][20] , \data_i[9][19] ,
         \data_i[9][18] , \data_i[9][17] , \data_i[9][16] , \data_i[9][15] ,
         \data_i[9][14] , \data_i[9][13] , \data_i[9][12] , \data_i[9][11] ,
         \data_i[9][10] , \data_i[9][9] , \data_i[9][8] , \data_i[9][7] ,
         \data_i[9][6] , \data_i[9][5] , \data_i[9][4] , \data_i[9][3] ,
         \data_i[9][2] , \data_i[9][1] , \data_i[9][0] , \data_i[8][31] ,
         \data_i[8][30] , \data_i[8][29] , \data_i[8][28] , \data_i[8][27] ,
         \data_i[8][26] , \data_i[8][25] , \data_i[8][24] , \data_i[8][23] ,
         \data_i[8][22] , \data_i[8][21] , \data_i[8][20] , \data_i[8][19] ,
         \data_i[8][18] , \data_i[8][17] , \data_i[8][16] , \data_i[8][15] ,
         \data_i[8][14] , \data_i[8][13] , \data_i[8][12] , \data_i[8][11] ,
         \data_i[8][10] , \data_i[8][9] , \data_i[8][8] , \data_i[8][7] ,
         \data_i[8][6] , \data_i[8][5] , \data_i[8][4] , \data_i[8][3] ,
         \data_i[8][2] , \data_i[8][1] , \data_i[8][0] , \data_i[7][31] ,
         \data_i[7][30] , \data_i[7][29] , \data_i[7][28] , \data_i[7][27] ,
         \data_i[7][26] , \data_i[7][25] , \data_i[7][24] , \data_i[7][23] ,
         \data_i[7][22] , \data_i[7][21] , \data_i[7][20] , \data_i[7][19] ,
         \data_i[7][18] , \data_i[7][17] , \data_i[7][16] , \data_i[7][15] ,
         \data_i[7][14] , \data_i[7][13] , \data_i[7][12] , \data_i[7][11] ,
         \data_i[7][10] , \data_i[7][9] , \data_i[7][8] , \data_i[7][7] ,
         \data_i[7][6] , \data_i[7][5] , \data_i[7][4] , \data_i[7][3] ,
         \data_i[7][2] , \data_i[7][1] , \data_i[7][0] , \data_i[6][31] ,
         \data_i[6][30] , \data_i[6][29] , \data_i[6][28] , \data_i[6][27] ,
         \data_i[6][26] , \data_i[6][25] , \data_i[6][24] , \data_i[6][23] ,
         \data_i[6][22] , \data_i[6][21] , \data_i[6][20] , \data_i[6][19] ,
         \data_i[6][18] , \data_i[6][17] , \data_i[6][16] , \data_i[6][15] ,
         \data_i[6][14] , \data_i[6][13] , \data_i[6][12] , \data_i[6][11] ,
         \data_i[6][10] , \data_i[6][9] , \data_i[6][8] , \data_i[6][7] ,
         \data_i[6][6] , \data_i[6][5] , \data_i[6][4] , \data_i[6][3] ,
         \data_i[6][2] , \data_i[6][1] , \data_i[6][0] , \data_i[5][31] ,
         \data_i[5][30] , \data_i[5][29] , \data_i[5][28] , \data_i[5][27] ,
         \data_i[5][26] , \data_i[5][25] , \data_i[5][24] , \data_i[5][23] ,
         \data_i[5][22] , \data_i[5][21] , \data_i[5][20] , \data_i[5][19] ,
         \data_i[5][18] , \data_i[5][17] , \data_i[5][16] , \data_i[5][15] ,
         \data_i[5][14] , \data_i[5][13] , \data_i[5][12] , \data_i[5][11] ,
         \data_i[5][10] , \data_i[5][9] , \data_i[5][8] , \data_i[5][7] ,
         \data_i[5][6] , \data_i[5][5] , \data_i[5][4] , \data_i[5][3] ,
         \data_i[5][2] , \data_i[5][1] , \data_i[5][0] , \data_i[4][31] ,
         \data_i[4][30] , \data_i[4][29] , \data_i[4][28] , \data_i[4][27] ,
         \data_i[4][26] , \data_i[4][25] , \data_i[4][24] , \data_i[4][23] ,
         \data_i[4][22] , \data_i[4][21] , \data_i[4][20] , \data_i[4][19] ,
         \data_i[4][18] , \data_i[4][17] , \data_i[4][16] , \data_i[4][15] ,
         \data_i[4][14] , \data_i[4][13] , \data_i[4][12] , \data_i[4][11] ,
         \data_i[4][10] , \data_i[4][9] , \data_i[4][8] , \data_i[4][7] ,
         \data_i[4][6] , \data_i[4][5] , \data_i[4][4] , \data_i[4][3] ,
         \data_i[4][2] , \data_i[4][1] , \data_i[4][0] , \data_i[3][31] ,
         \data_i[3][30] , \data_i[3][29] , \data_i[3][28] , \data_i[3][27] ,
         \data_i[3][26] , \data_i[3][25] , \data_i[3][24] , \data_i[3][23] ,
         \data_i[3][22] , \data_i[3][21] , \data_i[3][20] , \data_i[3][19] ,
         \data_i[3][18] , \data_i[3][17] , \data_i[3][16] , \data_i[3][15] ,
         \data_i[3][14] , \data_i[3][13] , \data_i[3][12] , \data_i[3][11] ,
         \data_i[3][10] , \data_i[3][9] , \data_i[3][8] , \data_i[3][7] ,
         \data_i[3][6] , \data_i[3][5] , \data_i[3][4] , \data_i[3][3] ,
         \data_i[3][2] , \data_i[3][1] , \data_i[3][0] , \data_i[2][31] ,
         \data_i[2][30] , \data_i[2][29] , \data_i[2][28] , \data_i[2][27] ,
         \data_i[2][26] , \data_i[2][25] , \data_i[2][24] , \data_i[2][23] ,
         \data_i[2][22] , \data_i[2][21] , \data_i[2][20] , \data_i[2][19] ,
         \data_i[2][18] , \data_i[2][17] , \data_i[2][16] , \data_i[2][15] ,
         \data_i[2][14] , \data_i[2][13] , \data_i[2][12] , \data_i[2][11] ,
         \data_i[2][10] , \data_i[2][9] , \data_i[2][8] , \data_i[2][7] ,
         \data_i[2][6] , \data_i[2][5] , \data_i[2][4] , \data_i[2][3] ,
         \data_i[2][2] , \data_i[2][1] , \data_i[2][0] , \data_i[1][31] ,
         \data_i[1][30] , \data_i[1][29] , \data_i[1][28] , \data_i[1][27] ,
         \data_i[1][26] , \data_i[1][25] , \data_i[1][24] , \data_i[1][23] ,
         \data_i[1][22] , \data_i[1][21] , \data_i[1][20] , \data_i[1][19] ,
         \data_i[1][18] , \data_i[1][17] , \data_i[1][16] , \data_i[1][15] ,
         \data_i[1][14] , \data_i[1][13] , \data_i[1][12] , \data_i[1][11] ,
         \data_i[1][10] , \data_i[1][9] , \data_i[1][8] , \data_i[1][7] ,
         \data_i[1][6] , \data_i[1][5] , \data_i[1][4] , \data_i[1][3] ,
         \data_i[1][2] , \data_i[1][1] , \data_i[1][0] , \data_i[0][31] ,
         \data_i[0][30] , \data_i[0][29] , \data_i[0][28] , \data_i[0][27] ,
         \data_i[0][26] , \data_i[0][25] , \data_i[0][24] , \data_i[0][23] ,
         \data_i[0][22] , \data_i[0][21] , \data_i[0][20] , \data_i[0][19] ,
         \data_i[0][18] , \data_i[0][17] , \data_i[0][16] , \data_i[0][15] ,
         \data_i[0][14] , \data_i[0][13] , \data_i[0][12] , \data_i[0][11] ,
         \data_i[0][10] , \data_i[0][9] , \data_i[0][8] , \data_i[0][7] ,
         \data_i[0][6] , \data_i[0][5] , \data_i[0][4] , \data_i[0][3] ,
         \data_i[0][2] , \data_i[0][1] , \data_i[0][0] ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690;

  NOR2X0 U1 ( .IN1(n42), .IN2(n50), .QN(n26) );
  NOR2X0 U2 ( .IN1(n49), .IN2(n42), .QN(n9) );
  NOR2X0 U3 ( .IN1(n43), .IN2(n49), .QN(n25) );
  NOR2X0 U4 ( .IN1(n42), .IN2(n51), .QN(n11) );
  NOR2X0 U5 ( .IN1(n43), .IN2(n51), .QN(n27) );
  NOR2X0 U6 ( .IN1(n43), .IN2(n50), .QN(n10) );
  NOR2X0 U7 ( .IN1(n42), .IN2(n52), .QN(n28) );
  NOR2X0 U8 ( .IN1(n49), .IN2(n60), .QN(n1) );
  NOR2X0 U9 ( .IN1(n42), .IN2(n58), .QN(n30) );
  NOR2X0 U10 ( .IN1(n42), .IN2(n57), .QN(n13) );
  NOR2X0 U11 ( .IN1(n50), .IN2(n60), .QN(n18) );
  NOR2X0 U12 ( .IN1(n59), .IN2(n60), .QN(n7) );
  NOR2X0 U13 ( .IN1(n43), .IN2(n57), .QN(n29) );
  NOR2X0 U14 ( .IN1(n42), .IN2(n59), .QN(n15) );
  NOR2X0 U15 ( .IN1(n57), .IN2(n60), .QN(n5) );
  NOR2X0 U16 ( .IN1(n50), .IN2(n61), .QN(n2) );
  NOR2X0 U17 ( .IN1(n57), .IN2(n61), .QN(n21) );
  NOR2X0 U18 ( .IN1(n62), .IN2(n60), .QN(n24) );
  NOR2X0 U19 ( .IN1(n49), .IN2(n61), .QN(n17) );
  NOR2X0 U20 ( .IN1(n43), .IN2(n59), .QN(n31) );
  NOR2X0 U21 ( .IN1(n43), .IN2(n58), .QN(n14) );
  NOR2X0 U22 ( .IN1(n58), .IN2(n61), .QN(n6) );
  NOR2X0 U23 ( .IN1(n62), .IN2(n61), .QN(n8) );
  NOR2X0 U24 ( .IN1(n58), .IN2(n60), .QN(n22) );
  NOR2X0 U25 ( .IN1(n52), .IN2(n61), .QN(n4) );
  NOR2X0 U26 ( .IN1(n43), .IN2(n62), .QN(n16) );
  NOR2X0 U27 ( .IN1(n42), .IN2(n62), .QN(n32) );
  NOR2X0 U28 ( .IN1(n43), .IN2(n52), .QN(n12) );
  NOR2X0 U29 ( .IN1(n51), .IN2(n61), .QN(n19) );
  NOR2X0 U30 ( .IN1(n59), .IN2(n61), .QN(n23) );
  NOR2X0 U31 ( .IN1(n52), .IN2(n60), .QN(n20) );
  NOR2X0 U32 ( .IN1(n51), .IN2(n60), .QN(n3) );
  INVX0 U33 ( .INP(select_i[2]), .ZN(n39) );
  INVX0 U34 ( .INP(select_i[0]), .ZN(n48) );
  INVX0 U35 ( .INP(select_i[4]), .ZN(n33) );
  NAND2X1 U36 ( .IN1(select_i[4]), .IN2(n48), .QN(n61) );
  NAND2X1 U37 ( .IN1(select_i[2]), .IN2(n41), .QN(n62) );
  NAND2X1 U38 ( .IN1(n41), .IN2(n39), .QN(n58) );
  NAND2X1 U39 ( .IN1(select_i[0]), .IN2(n33), .QN(n42) );
  NAND2X1 U40 ( .IN1(n33), .IN2(n48), .QN(n43) );
  NAND2X1 U41 ( .IN1(select_i[4]), .IN2(select_i[0]), .QN(n60) );
  NAND3X0 U42 ( .IN1(select_i[1]), .IN2(select_i[3]), .IN3(n39), .QN(n49) );
  AO22X1 U43 ( .IN1(n25), .IN2(\data_i[10][0] ), .IN3(n9), .IN4(
        \data_i[11][0] ), .Q(n38) );
  INVX0 U44 ( .INP(select_i[1]), .ZN(n34) );
  NAND3X0 U45 ( .IN1(select_i[3]), .IN2(n39), .IN3(n34), .QN(n50) );
  AO22X1 U46 ( .IN1(n26), .IN2(\data_i[9][0] ), .IN3(n10), .IN4(\data_i[8][0] ), .Q(n37) );
  NAND3X0 U47 ( .IN1(select_i[2]), .IN2(select_i[1]), .IN3(select_i[3]), .QN(
        n51) );
  AO22X1 U48 ( .IN1(n27), .IN2(\data_i[14][0] ), .IN3(n11), .IN4(
        \data_i[15][0] ), .Q(n36) );
  NAND3X0 U49 ( .IN1(select_i[2]), .IN2(select_i[3]), .IN3(n34), .QN(n52) );
  AO22X1 U50 ( .IN1(n28), .IN2(\data_i[13][0] ), .IN3(n12), .IN4(
        \data_i[12][0] ), .Q(n35) );
  NOR4X0 U51 ( .IN1(n38), .IN2(n37), .IN3(n36), .IN4(n35), .QN(n70) );
  INVX0 U52 ( .INP(select_i[3]), .ZN(n40) );
  NAND3X0 U53 ( .IN1(select_i[1]), .IN2(n39), .IN3(n40), .QN(n57) );
  AO22X1 U54 ( .IN1(n29), .IN2(\data_i[2][0] ), .IN3(n13), .IN4(\data_i[3][0] ), .Q(n47) );
  NOR2X0 U55 ( .IN1(select_i[1]), .IN2(select_i[3]), .QN(n41) );
  AO22X1 U56 ( .IN1(n30), .IN2(\data_i[1][0] ), .IN3(n14), .IN4(\data_i[0][0] ), .Q(n46) );
  NAND3X0 U57 ( .IN1(select_i[1]), .IN2(select_i[2]), .IN3(n40), .QN(n59) );
  AO22X1 U58 ( .IN1(n31), .IN2(\data_i[6][0] ), .IN3(n15), .IN4(\data_i[7][0] ), .Q(n45) );
  AO22X1 U59 ( .IN1(n32), .IN2(\data_i[5][0] ), .IN3(n16), .IN4(\data_i[4][0] ), .Q(n44) );
  NOR4X0 U60 ( .IN1(n47), .IN2(n46), .IN3(n45), .IN4(n44), .QN(n69) );
  AO22X1 U61 ( .IN1(n17), .IN2(\data_i[26][0] ), .IN3(n1), .IN4(
        \data_i[27][0] ), .Q(n56) );
  AO22X1 U62 ( .IN1(n18), .IN2(\data_i[25][0] ), .IN3(n2), .IN4(
        \data_i[24][0] ), .Q(n55) );
  AO22X1 U63 ( .IN1(n19), .IN2(\data_i[30][0] ), .IN3(n3), .IN4(
        \data_i[31][0] ), .Q(n54) );
  AO22X1 U64 ( .IN1(n20), .IN2(\data_i[29][0] ), .IN3(n4), .IN4(
        \data_i[28][0] ), .Q(n53) );
  NOR4X0 U65 ( .IN1(n56), .IN2(n55), .IN3(n54), .IN4(n53), .QN(n68) );
  AO22X1 U66 ( .IN1(n21), .IN2(\data_i[18][0] ), .IN3(n5), .IN4(
        \data_i[19][0] ), .Q(n66) );
  AO22X1 U67 ( .IN1(n22), .IN2(\data_i[17][0] ), .IN3(n6), .IN4(
        \data_i[16][0] ), .Q(n65) );
  AO22X1 U68 ( .IN1(n23), .IN2(\data_i[22][0] ), .IN3(n7), .IN4(
        \data_i[23][0] ), .Q(n64) );
  AO22X1 U69 ( .IN1(n24), .IN2(\data_i[21][0] ), .IN3(n8), .IN4(
        \data_i[20][0] ), .Q(n63) );
  NOR4X0 U70 ( .IN1(n66), .IN2(n65), .IN3(n64), .IN4(n63), .QN(n67) );
  NAND4X0 U71 ( .IN1(n70), .IN2(n69), .IN3(n68), .IN4(n67), .QN(data_o[0]) );
  AO22X1 U72 ( .IN1(n25), .IN2(\data_i[10][10] ), .IN3(n9), .IN4(
        \data_i[11][10] ), .Q(n74) );
  AO22X1 U73 ( .IN1(n26), .IN2(\data_i[9][10] ), .IN3(n10), .IN4(
        \data_i[8][10] ), .Q(n73) );
  AO22X1 U74 ( .IN1(n27), .IN2(\data_i[14][10] ), .IN3(n11), .IN4(
        \data_i[15][10] ), .Q(n72) );
  AO22X1 U75 ( .IN1(n28), .IN2(\data_i[13][10] ), .IN3(n12), .IN4(
        \data_i[12][10] ), .Q(n71) );
  NOR4X0 U76 ( .IN1(n74), .IN2(n73), .IN3(n72), .IN4(n71), .QN(n90) );
  AO22X1 U77 ( .IN1(n29), .IN2(\data_i[2][10] ), .IN3(n13), .IN4(
        \data_i[3][10] ), .Q(n78) );
  AO22X1 U78 ( .IN1(n30), .IN2(\data_i[1][10] ), .IN3(n14), .IN4(
        \data_i[0][10] ), .Q(n77) );
  AO22X1 U79 ( .IN1(n31), .IN2(\data_i[6][10] ), .IN3(n15), .IN4(
        \data_i[7][10] ), .Q(n76) );
  AO22X1 U80 ( .IN1(n32), .IN2(\data_i[5][10] ), .IN3(n16), .IN4(
        \data_i[4][10] ), .Q(n75) );
  NOR4X0 U81 ( .IN1(n78), .IN2(n77), .IN3(n76), .IN4(n75), .QN(n89) );
  AO22X1 U82 ( .IN1(n17), .IN2(\data_i[26][10] ), .IN3(n1), .IN4(
        \data_i[27][10] ), .Q(n82) );
  AO22X1 U83 ( .IN1(n18), .IN2(\data_i[25][10] ), .IN3(n2), .IN4(
        \data_i[24][10] ), .Q(n81) );
  AO22X1 U84 ( .IN1(n19), .IN2(\data_i[30][10] ), .IN3(n3), .IN4(
        \data_i[31][10] ), .Q(n80) );
  AO22X1 U85 ( .IN1(n20), .IN2(\data_i[29][10] ), .IN3(n4), .IN4(
        \data_i[28][10] ), .Q(n79) );
  NOR4X0 U86 ( .IN1(n82), .IN2(n81), .IN3(n80), .IN4(n79), .QN(n88) );
  AO22X1 U87 ( .IN1(n21), .IN2(\data_i[18][10] ), .IN3(n5), .IN4(
        \data_i[19][10] ), .Q(n86) );
  AO22X1 U88 ( .IN1(n22), .IN2(\data_i[17][10] ), .IN3(n6), .IN4(
        \data_i[16][10] ), .Q(n85) );
  AO22X1 U89 ( .IN1(n23), .IN2(\data_i[22][10] ), .IN3(n7), .IN4(
        \data_i[23][10] ), .Q(n84) );
  AO22X1 U90 ( .IN1(n24), .IN2(\data_i[21][10] ), .IN3(n8), .IN4(
        \data_i[20][10] ), .Q(n83) );
  NOR4X0 U91 ( .IN1(n86), .IN2(n85), .IN3(n84), .IN4(n83), .QN(n87) );
  NAND4X0 U92 ( .IN1(n90), .IN2(n89), .IN3(n88), .IN4(n87), .QN(data_o[10]) );
  AO22X1 U93 ( .IN1(n25), .IN2(\data_i[10][11] ), .IN3(n9), .IN4(
        \data_i[11][11] ), .Q(n94) );
  AO22X1 U94 ( .IN1(n26), .IN2(\data_i[9][11] ), .IN3(n10), .IN4(
        \data_i[8][11] ), .Q(n93) );
  AO22X1 U95 ( .IN1(n27), .IN2(\data_i[14][11] ), .IN3(n11), .IN4(
        \data_i[15][11] ), .Q(n92) );
  AO22X1 U96 ( .IN1(n28), .IN2(\data_i[13][11] ), .IN3(n12), .IN4(
        \data_i[12][11] ), .Q(n91) );
  NOR4X0 U97 ( .IN1(n94), .IN2(n93), .IN3(n92), .IN4(n91), .QN(n110) );
  AO22X1 U98 ( .IN1(n29), .IN2(\data_i[2][11] ), .IN3(n13), .IN4(
        \data_i[3][11] ), .Q(n98) );
  AO22X1 U99 ( .IN1(n30), .IN2(\data_i[1][11] ), .IN3(n14), .IN4(
        \data_i[0][11] ), .Q(n97) );
  AO22X1 U100 ( .IN1(n31), .IN2(\data_i[6][11] ), .IN3(n15), .IN4(
        \data_i[7][11] ), .Q(n96) );
  AO22X1 U101 ( .IN1(n32), .IN2(\data_i[5][11] ), .IN3(n16), .IN4(
        \data_i[4][11] ), .Q(n95) );
  NOR4X0 U102 ( .IN1(n98), .IN2(n97), .IN3(n96), .IN4(n95), .QN(n109) );
  AO22X1 U103 ( .IN1(n17), .IN2(\data_i[26][11] ), .IN3(n1), .IN4(
        \data_i[27][11] ), .Q(n102) );
  AO22X1 U104 ( .IN1(n18), .IN2(\data_i[25][11] ), .IN3(n2), .IN4(
        \data_i[24][11] ), .Q(n101) );
  AO22X1 U105 ( .IN1(n19), .IN2(\data_i[30][11] ), .IN3(n3), .IN4(
        \data_i[31][11] ), .Q(n100) );
  AO22X1 U106 ( .IN1(n20), .IN2(\data_i[29][11] ), .IN3(n4), .IN4(
        \data_i[28][11] ), .Q(n99) );
  NOR4X0 U107 ( .IN1(n102), .IN2(n101), .IN3(n100), .IN4(n99), .QN(n108) );
  AO22X1 U108 ( .IN1(n21), .IN2(\data_i[18][11] ), .IN3(n5), .IN4(
        \data_i[19][11] ), .Q(n106) );
  AO22X1 U109 ( .IN1(n22), .IN2(\data_i[17][11] ), .IN3(n6), .IN4(
        \data_i[16][11] ), .Q(n105) );
  AO22X1 U110 ( .IN1(n23), .IN2(\data_i[22][11] ), .IN3(n7), .IN4(
        \data_i[23][11] ), .Q(n104) );
  AO22X1 U111 ( .IN1(n24), .IN2(\data_i[21][11] ), .IN3(n8), .IN4(
        \data_i[20][11] ), .Q(n103) );
  NOR4X0 U112 ( .IN1(n106), .IN2(n105), .IN3(n104), .IN4(n103), .QN(n107) );
  NAND4X0 U113 ( .IN1(n110), .IN2(n109), .IN3(n108), .IN4(n107), .QN(
        data_o[11]) );
  AO22X1 U114 ( .IN1(n25), .IN2(\data_i[10][12] ), .IN3(n9), .IN4(
        \data_i[11][12] ), .Q(n114) );
  AO22X1 U115 ( .IN1(n26), .IN2(\data_i[9][12] ), .IN3(n10), .IN4(
        \data_i[8][12] ), .Q(n113) );
  AO22X1 U116 ( .IN1(n27), .IN2(\data_i[14][12] ), .IN3(n11), .IN4(
        \data_i[15][12] ), .Q(n112) );
  AO22X1 U117 ( .IN1(n28), .IN2(\data_i[13][12] ), .IN3(n12), .IN4(
        \data_i[12][12] ), .Q(n111) );
  NOR4X0 U118 ( .IN1(n114), .IN2(n113), .IN3(n112), .IN4(n111), .QN(n130) );
  AO22X1 U119 ( .IN1(n29), .IN2(\data_i[2][12] ), .IN3(n13), .IN4(
        \data_i[3][12] ), .Q(n118) );
  AO22X1 U120 ( .IN1(n30), .IN2(\data_i[1][12] ), .IN3(n14), .IN4(
        \data_i[0][12] ), .Q(n117) );
  AO22X1 U121 ( .IN1(n31), .IN2(\data_i[6][12] ), .IN3(n15), .IN4(
        \data_i[7][12] ), .Q(n116) );
  AO22X1 U122 ( .IN1(n32), .IN2(\data_i[5][12] ), .IN3(n16), .IN4(
        \data_i[4][12] ), .Q(n115) );
  NOR4X0 U123 ( .IN1(n118), .IN2(n117), .IN3(n116), .IN4(n115), .QN(n129) );
  AO22X1 U124 ( .IN1(n17), .IN2(\data_i[26][12] ), .IN3(n1), .IN4(
        \data_i[27][12] ), .Q(n122) );
  AO22X1 U125 ( .IN1(n18), .IN2(\data_i[25][12] ), .IN3(n2), .IN4(
        \data_i[24][12] ), .Q(n121) );
  AO22X1 U126 ( .IN1(n19), .IN2(\data_i[30][12] ), .IN3(n3), .IN4(
        \data_i[31][12] ), .Q(n120) );
  AO22X1 U127 ( .IN1(n20), .IN2(\data_i[29][12] ), .IN3(n4), .IN4(
        \data_i[28][12] ), .Q(n119) );
  NOR4X0 U128 ( .IN1(n122), .IN2(n121), .IN3(n120), .IN4(n119), .QN(n128) );
  AO22X1 U129 ( .IN1(n21), .IN2(\data_i[18][12] ), .IN3(n5), .IN4(
        \data_i[19][12] ), .Q(n126) );
  AO22X1 U130 ( .IN1(n22), .IN2(\data_i[17][12] ), .IN3(n6), .IN4(
        \data_i[16][12] ), .Q(n125) );
  AO22X1 U131 ( .IN1(n23), .IN2(\data_i[22][12] ), .IN3(n7), .IN4(
        \data_i[23][12] ), .Q(n124) );
  AO22X1 U132 ( .IN1(n24), .IN2(\data_i[21][12] ), .IN3(n8), .IN4(
        \data_i[20][12] ), .Q(n123) );
  NOR4X0 U133 ( .IN1(n126), .IN2(n125), .IN3(n124), .IN4(n123), .QN(n127) );
  NAND4X0 U134 ( .IN1(n130), .IN2(n129), .IN3(n128), .IN4(n127), .QN(
        data_o[12]) );
  AO22X1 U135 ( .IN1(n25), .IN2(\data_i[10][13] ), .IN3(n9), .IN4(
        \data_i[11][13] ), .Q(n134) );
  AO22X1 U136 ( .IN1(n26), .IN2(\data_i[9][13] ), .IN3(n10), .IN4(
        \data_i[8][13] ), .Q(n133) );
  AO22X1 U137 ( .IN1(n27), .IN2(\data_i[14][13] ), .IN3(n11), .IN4(
        \data_i[15][13] ), .Q(n132) );
  AO22X1 U138 ( .IN1(n28), .IN2(\data_i[13][13] ), .IN3(n12), .IN4(
        \data_i[12][13] ), .Q(n131) );
  NOR4X0 U139 ( .IN1(n134), .IN2(n133), .IN3(n132), .IN4(n131), .QN(n150) );
  AO22X1 U140 ( .IN1(n29), .IN2(\data_i[2][13] ), .IN3(n13), .IN4(
        \data_i[3][13] ), .Q(n138) );
  AO22X1 U141 ( .IN1(n30), .IN2(\data_i[1][13] ), .IN3(n14), .IN4(
        \data_i[0][13] ), .Q(n137) );
  AO22X1 U142 ( .IN1(n31), .IN2(\data_i[6][13] ), .IN3(n15), .IN4(
        \data_i[7][13] ), .Q(n136) );
  AO22X1 U143 ( .IN1(n32), .IN2(\data_i[5][13] ), .IN3(n16), .IN4(
        \data_i[4][13] ), .Q(n135) );
  NOR4X0 U144 ( .IN1(n138), .IN2(n137), .IN3(n136), .IN4(n135), .QN(n149) );
  AO22X1 U145 ( .IN1(n17), .IN2(\data_i[26][13] ), .IN3(n1), .IN4(
        \data_i[27][13] ), .Q(n142) );
  AO22X1 U146 ( .IN1(n18), .IN2(\data_i[25][13] ), .IN3(n2), .IN4(
        \data_i[24][13] ), .Q(n141) );
  AO22X1 U147 ( .IN1(n19), .IN2(\data_i[30][13] ), .IN3(n3), .IN4(
        \data_i[31][13] ), .Q(n140) );
  AO22X1 U148 ( .IN1(n20), .IN2(\data_i[29][13] ), .IN3(n4), .IN4(
        \data_i[28][13] ), .Q(n139) );
  NOR4X0 U149 ( .IN1(n142), .IN2(n141), .IN3(n140), .IN4(n139), .QN(n148) );
  AO22X1 U150 ( .IN1(n21), .IN2(\data_i[18][13] ), .IN3(n5), .IN4(
        \data_i[19][13] ), .Q(n146) );
  AO22X1 U151 ( .IN1(n22), .IN2(\data_i[17][13] ), .IN3(n6), .IN4(
        \data_i[16][13] ), .Q(n145) );
  AO22X1 U152 ( .IN1(n23), .IN2(\data_i[22][13] ), .IN3(n7), .IN4(
        \data_i[23][13] ), .Q(n144) );
  AO22X1 U153 ( .IN1(n24), .IN2(\data_i[21][13] ), .IN3(n8), .IN4(
        \data_i[20][13] ), .Q(n143) );
  NOR4X0 U154 ( .IN1(n146), .IN2(n145), .IN3(n144), .IN4(n143), .QN(n147) );
  NAND4X0 U155 ( .IN1(n150), .IN2(n149), .IN3(n148), .IN4(n147), .QN(
        data_o[13]) );
  AO22X1 U156 ( .IN1(n25), .IN2(\data_i[10][14] ), .IN3(n9), .IN4(
        \data_i[11][14] ), .Q(n154) );
  AO22X1 U157 ( .IN1(n26), .IN2(\data_i[9][14] ), .IN3(n10), .IN4(
        \data_i[8][14] ), .Q(n153) );
  AO22X1 U158 ( .IN1(n27), .IN2(\data_i[14][14] ), .IN3(n11), .IN4(
        \data_i[15][14] ), .Q(n152) );
  AO22X1 U159 ( .IN1(n28), .IN2(\data_i[13][14] ), .IN3(n12), .IN4(
        \data_i[12][14] ), .Q(n151) );
  NOR4X0 U160 ( .IN1(n154), .IN2(n153), .IN3(n152), .IN4(n151), .QN(n170) );
  AO22X1 U161 ( .IN1(n29), .IN2(\data_i[2][14] ), .IN3(n13), .IN4(
        \data_i[3][14] ), .Q(n158) );
  AO22X1 U162 ( .IN1(n30), .IN2(\data_i[1][14] ), .IN3(n14), .IN4(
        \data_i[0][14] ), .Q(n157) );
  AO22X1 U163 ( .IN1(n31), .IN2(\data_i[6][14] ), .IN3(n15), .IN4(
        \data_i[7][14] ), .Q(n156) );
  AO22X1 U164 ( .IN1(n32), .IN2(\data_i[5][14] ), .IN3(n16), .IN4(
        \data_i[4][14] ), .Q(n155) );
  NOR4X0 U165 ( .IN1(n158), .IN2(n157), .IN3(n156), .IN4(n155), .QN(n169) );
  AO22X1 U166 ( .IN1(n17), .IN2(\data_i[26][14] ), .IN3(n1), .IN4(
        \data_i[27][14] ), .Q(n162) );
  AO22X1 U167 ( .IN1(n18), .IN2(\data_i[25][14] ), .IN3(n2), .IN4(
        \data_i[24][14] ), .Q(n161) );
  AO22X1 U168 ( .IN1(n19), .IN2(\data_i[30][14] ), .IN3(n3), .IN4(
        \data_i[31][14] ), .Q(n160) );
  AO22X1 U169 ( .IN1(n20), .IN2(\data_i[29][14] ), .IN3(n4), .IN4(
        \data_i[28][14] ), .Q(n159) );
  NOR4X0 U170 ( .IN1(n162), .IN2(n161), .IN3(n160), .IN4(n159), .QN(n168) );
  AO22X1 U171 ( .IN1(n21), .IN2(\data_i[18][14] ), .IN3(n5), .IN4(
        \data_i[19][14] ), .Q(n166) );
  AO22X1 U172 ( .IN1(n22), .IN2(\data_i[17][14] ), .IN3(n6), .IN4(
        \data_i[16][14] ), .Q(n165) );
  AO22X1 U173 ( .IN1(n23), .IN2(\data_i[22][14] ), .IN3(n7), .IN4(
        \data_i[23][14] ), .Q(n164) );
  AO22X1 U174 ( .IN1(n24), .IN2(\data_i[21][14] ), .IN3(n8), .IN4(
        \data_i[20][14] ), .Q(n163) );
  NOR4X0 U175 ( .IN1(n166), .IN2(n165), .IN3(n164), .IN4(n163), .QN(n167) );
  NAND4X0 U176 ( .IN1(n170), .IN2(n169), .IN3(n168), .IN4(n167), .QN(
        data_o[14]) );
  AO22X1 U177 ( .IN1(n25), .IN2(\data_i[10][15] ), .IN3(n9), .IN4(
        \data_i[11][15] ), .Q(n174) );
  AO22X1 U178 ( .IN1(n26), .IN2(\data_i[9][15] ), .IN3(n10), .IN4(
        \data_i[8][15] ), .Q(n173) );
  AO22X1 U179 ( .IN1(n27), .IN2(\data_i[14][15] ), .IN3(n11), .IN4(
        \data_i[15][15] ), .Q(n172) );
  AO22X1 U180 ( .IN1(n28), .IN2(\data_i[13][15] ), .IN3(n12), .IN4(
        \data_i[12][15] ), .Q(n171) );
  NOR4X0 U181 ( .IN1(n174), .IN2(n173), .IN3(n172), .IN4(n171), .QN(n190) );
  AO22X1 U182 ( .IN1(n29), .IN2(\data_i[2][15] ), .IN3(n13), .IN4(
        \data_i[3][15] ), .Q(n178) );
  AO22X1 U183 ( .IN1(n30), .IN2(\data_i[1][15] ), .IN3(n14), .IN4(
        \data_i[0][15] ), .Q(n177) );
  AO22X1 U184 ( .IN1(n31), .IN2(\data_i[6][15] ), .IN3(n15), .IN4(
        \data_i[7][15] ), .Q(n176) );
  AO22X1 U185 ( .IN1(n32), .IN2(\data_i[5][15] ), .IN3(n16), .IN4(
        \data_i[4][15] ), .Q(n175) );
  NOR4X0 U186 ( .IN1(n178), .IN2(n177), .IN3(n176), .IN4(n175), .QN(n189) );
  AO22X1 U187 ( .IN1(n17), .IN2(\data_i[26][15] ), .IN3(n1), .IN4(
        \data_i[27][15] ), .Q(n182) );
  AO22X1 U188 ( .IN1(n18), .IN2(\data_i[25][15] ), .IN3(n2), .IN4(
        \data_i[24][15] ), .Q(n181) );
  AO22X1 U189 ( .IN1(n19), .IN2(\data_i[30][15] ), .IN3(n3), .IN4(
        \data_i[31][15] ), .Q(n180) );
  AO22X1 U190 ( .IN1(n20), .IN2(\data_i[29][15] ), .IN3(n4), .IN4(
        \data_i[28][15] ), .Q(n179) );
  NOR4X0 U191 ( .IN1(n182), .IN2(n181), .IN3(n180), .IN4(n179), .QN(n188) );
  AO22X1 U192 ( .IN1(n21), .IN2(\data_i[18][15] ), .IN3(n5), .IN4(
        \data_i[19][15] ), .Q(n186) );
  AO22X1 U193 ( .IN1(n22), .IN2(\data_i[17][15] ), .IN3(n6), .IN4(
        \data_i[16][15] ), .Q(n185) );
  AO22X1 U194 ( .IN1(n23), .IN2(\data_i[22][15] ), .IN3(n7), .IN4(
        \data_i[23][15] ), .Q(n184) );
  AO22X1 U195 ( .IN1(n24), .IN2(\data_i[21][15] ), .IN3(n8), .IN4(
        \data_i[20][15] ), .Q(n183) );
  NOR4X0 U196 ( .IN1(n186), .IN2(n185), .IN3(n184), .IN4(n183), .QN(n187) );
  NAND4X0 U197 ( .IN1(n190), .IN2(n189), .IN3(n188), .IN4(n187), .QN(
        data_o[15]) );
  AO22X1 U198 ( .IN1(n25), .IN2(\data_i[10][16] ), .IN3(n9), .IN4(
        \data_i[11][16] ), .Q(n194) );
  AO22X1 U199 ( .IN1(n26), .IN2(\data_i[9][16] ), .IN3(n10), .IN4(
        \data_i[8][16] ), .Q(n193) );
  AO22X1 U200 ( .IN1(n27), .IN2(\data_i[14][16] ), .IN3(n11), .IN4(
        \data_i[15][16] ), .Q(n192) );
  AO22X1 U201 ( .IN1(n28), .IN2(\data_i[13][16] ), .IN3(n12), .IN4(
        \data_i[12][16] ), .Q(n191) );
  NOR4X0 U202 ( .IN1(n194), .IN2(n193), .IN3(n192), .IN4(n191), .QN(n210) );
  AO22X1 U203 ( .IN1(n29), .IN2(\data_i[2][16] ), .IN3(n13), .IN4(
        \data_i[3][16] ), .Q(n198) );
  AO22X1 U204 ( .IN1(n30), .IN2(\data_i[1][16] ), .IN3(n14), .IN4(
        \data_i[0][16] ), .Q(n197) );
  AO22X1 U205 ( .IN1(n31), .IN2(\data_i[6][16] ), .IN3(n15), .IN4(
        \data_i[7][16] ), .Q(n196) );
  AO22X1 U206 ( .IN1(n32), .IN2(\data_i[5][16] ), .IN3(n16), .IN4(
        \data_i[4][16] ), .Q(n195) );
  NOR4X0 U207 ( .IN1(n198), .IN2(n197), .IN3(n196), .IN4(n195), .QN(n209) );
  AO22X1 U208 ( .IN1(n17), .IN2(\data_i[26][16] ), .IN3(n1), .IN4(
        \data_i[27][16] ), .Q(n202) );
  AO22X1 U209 ( .IN1(n18), .IN2(\data_i[25][16] ), .IN3(n2), .IN4(
        \data_i[24][16] ), .Q(n201) );
  AO22X1 U210 ( .IN1(n19), .IN2(\data_i[30][16] ), .IN3(n3), .IN4(
        \data_i[31][16] ), .Q(n200) );
  AO22X1 U211 ( .IN1(n20), .IN2(\data_i[29][16] ), .IN3(n4), .IN4(
        \data_i[28][16] ), .Q(n199) );
  NOR4X0 U212 ( .IN1(n202), .IN2(n201), .IN3(n200), .IN4(n199), .QN(n208) );
  AO22X1 U213 ( .IN1(n21), .IN2(\data_i[18][16] ), .IN3(n5), .IN4(
        \data_i[19][16] ), .Q(n206) );
  AO22X1 U214 ( .IN1(n22), .IN2(\data_i[17][16] ), .IN3(n6), .IN4(
        \data_i[16][16] ), .Q(n205) );
  AO22X1 U215 ( .IN1(n23), .IN2(\data_i[22][16] ), .IN3(n7), .IN4(
        \data_i[23][16] ), .Q(n204) );
  AO22X1 U216 ( .IN1(n24), .IN2(\data_i[21][16] ), .IN3(n8), .IN4(
        \data_i[20][16] ), .Q(n203) );
  NOR4X0 U217 ( .IN1(n206), .IN2(n205), .IN3(n204), .IN4(n203), .QN(n207) );
  NAND4X0 U218 ( .IN1(n210), .IN2(n209), .IN3(n208), .IN4(n207), .QN(
        data_o[16]) );
  AO22X1 U219 ( .IN1(n25), .IN2(\data_i[10][17] ), .IN3(n9), .IN4(
        \data_i[11][17] ), .Q(n214) );
  AO22X1 U220 ( .IN1(n26), .IN2(\data_i[9][17] ), .IN3(n10), .IN4(
        \data_i[8][17] ), .Q(n213) );
  AO22X1 U221 ( .IN1(n27), .IN2(\data_i[14][17] ), .IN3(n11), .IN4(
        \data_i[15][17] ), .Q(n212) );
  AO22X1 U222 ( .IN1(n28), .IN2(\data_i[13][17] ), .IN3(n12), .IN4(
        \data_i[12][17] ), .Q(n211) );
  NOR4X0 U223 ( .IN1(n214), .IN2(n213), .IN3(n212), .IN4(n211), .QN(n230) );
  AO22X1 U224 ( .IN1(n29), .IN2(\data_i[2][17] ), .IN3(n13), .IN4(
        \data_i[3][17] ), .Q(n218) );
  AO22X1 U225 ( .IN1(n30), .IN2(\data_i[1][17] ), .IN3(n14), .IN4(
        \data_i[0][17] ), .Q(n217) );
  AO22X1 U226 ( .IN1(n31), .IN2(\data_i[6][17] ), .IN3(n15), .IN4(
        \data_i[7][17] ), .Q(n216) );
  AO22X1 U227 ( .IN1(n32), .IN2(\data_i[5][17] ), .IN3(n16), .IN4(
        \data_i[4][17] ), .Q(n215) );
  NOR4X0 U228 ( .IN1(n218), .IN2(n217), .IN3(n216), .IN4(n215), .QN(n229) );
  AO22X1 U229 ( .IN1(n17), .IN2(\data_i[26][17] ), .IN3(n1), .IN4(
        \data_i[27][17] ), .Q(n222) );
  AO22X1 U230 ( .IN1(n18), .IN2(\data_i[25][17] ), .IN3(n2), .IN4(
        \data_i[24][17] ), .Q(n221) );
  AO22X1 U231 ( .IN1(n19), .IN2(\data_i[30][17] ), .IN3(n3), .IN4(
        \data_i[31][17] ), .Q(n220) );
  AO22X1 U232 ( .IN1(n20), .IN2(\data_i[29][17] ), .IN3(n4), .IN4(
        \data_i[28][17] ), .Q(n219) );
  NOR4X0 U233 ( .IN1(n222), .IN2(n221), .IN3(n220), .IN4(n219), .QN(n228) );
  AO22X1 U234 ( .IN1(n21), .IN2(\data_i[18][17] ), .IN3(n5), .IN4(
        \data_i[19][17] ), .Q(n226) );
  AO22X1 U235 ( .IN1(n22), .IN2(\data_i[17][17] ), .IN3(n6), .IN4(
        \data_i[16][17] ), .Q(n225) );
  AO22X1 U236 ( .IN1(n23), .IN2(\data_i[22][17] ), .IN3(n7), .IN4(
        \data_i[23][17] ), .Q(n224) );
  AO22X1 U237 ( .IN1(n24), .IN2(\data_i[21][17] ), .IN3(n8), .IN4(
        \data_i[20][17] ), .Q(n223) );
  NOR4X0 U238 ( .IN1(n226), .IN2(n225), .IN3(n224), .IN4(n223), .QN(n227) );
  NAND4X0 U239 ( .IN1(n230), .IN2(n229), .IN3(n228), .IN4(n227), .QN(
        data_o[17]) );
  AO22X1 U240 ( .IN1(n25), .IN2(\data_i[10][18] ), .IN3(n9), .IN4(
        \data_i[11][18] ), .Q(n234) );
  AO22X1 U241 ( .IN1(n26), .IN2(\data_i[9][18] ), .IN3(n10), .IN4(
        \data_i[8][18] ), .Q(n233) );
  AO22X1 U242 ( .IN1(n27), .IN2(\data_i[14][18] ), .IN3(n11), .IN4(
        \data_i[15][18] ), .Q(n232) );
  AO22X1 U243 ( .IN1(n28), .IN2(\data_i[13][18] ), .IN3(n12), .IN4(
        \data_i[12][18] ), .Q(n231) );
  NOR4X0 U244 ( .IN1(n234), .IN2(n233), .IN3(n232), .IN4(n231), .QN(n250) );
  AO22X1 U245 ( .IN1(n29), .IN2(\data_i[2][18] ), .IN3(n13), .IN4(
        \data_i[3][18] ), .Q(n238) );
  AO22X1 U246 ( .IN1(n30), .IN2(\data_i[1][18] ), .IN3(n14), .IN4(
        \data_i[0][18] ), .Q(n237) );
  AO22X1 U247 ( .IN1(n31), .IN2(\data_i[6][18] ), .IN3(n15), .IN4(
        \data_i[7][18] ), .Q(n236) );
  AO22X1 U248 ( .IN1(n32), .IN2(\data_i[5][18] ), .IN3(n16), .IN4(
        \data_i[4][18] ), .Q(n235) );
  NOR4X0 U249 ( .IN1(n238), .IN2(n237), .IN3(n236), .IN4(n235), .QN(n249) );
  AO22X1 U250 ( .IN1(n17), .IN2(\data_i[26][18] ), .IN3(n1), .IN4(
        \data_i[27][18] ), .Q(n242) );
  AO22X1 U251 ( .IN1(n18), .IN2(\data_i[25][18] ), .IN3(n2), .IN4(
        \data_i[24][18] ), .Q(n241) );
  AO22X1 U252 ( .IN1(n19), .IN2(\data_i[30][18] ), .IN3(n3), .IN4(
        \data_i[31][18] ), .Q(n240) );
  AO22X1 U253 ( .IN1(n20), .IN2(\data_i[29][18] ), .IN3(n4), .IN4(
        \data_i[28][18] ), .Q(n239) );
  NOR4X0 U254 ( .IN1(n242), .IN2(n241), .IN3(n240), .IN4(n239), .QN(n248) );
  AO22X1 U255 ( .IN1(n21), .IN2(\data_i[18][18] ), .IN3(n5), .IN4(
        \data_i[19][18] ), .Q(n246) );
  AO22X1 U256 ( .IN1(n22), .IN2(\data_i[17][18] ), .IN3(n6), .IN4(
        \data_i[16][18] ), .Q(n245) );
  AO22X1 U257 ( .IN1(n23), .IN2(\data_i[22][18] ), .IN3(n7), .IN4(
        \data_i[23][18] ), .Q(n244) );
  AO22X1 U258 ( .IN1(n24), .IN2(\data_i[21][18] ), .IN3(n8), .IN4(
        \data_i[20][18] ), .Q(n243) );
  NOR4X0 U259 ( .IN1(n246), .IN2(n245), .IN3(n244), .IN4(n243), .QN(n247) );
  NAND4X0 U260 ( .IN1(n250), .IN2(n249), .IN3(n248), .IN4(n247), .QN(
        data_o[18]) );
  AO22X1 U261 ( .IN1(n25), .IN2(\data_i[10][19] ), .IN3(n9), .IN4(
        \data_i[11][19] ), .Q(n254) );
  AO22X1 U262 ( .IN1(n26), .IN2(\data_i[9][19] ), .IN3(n10), .IN4(
        \data_i[8][19] ), .Q(n253) );
  AO22X1 U263 ( .IN1(n27), .IN2(\data_i[14][19] ), .IN3(n11), .IN4(
        \data_i[15][19] ), .Q(n252) );
  AO22X1 U264 ( .IN1(n28), .IN2(\data_i[13][19] ), .IN3(n12), .IN4(
        \data_i[12][19] ), .Q(n251) );
  NOR4X0 U265 ( .IN1(n254), .IN2(n253), .IN3(n252), .IN4(n251), .QN(n270) );
  AO22X1 U266 ( .IN1(n29), .IN2(\data_i[2][19] ), .IN3(n13), .IN4(
        \data_i[3][19] ), .Q(n258) );
  AO22X1 U267 ( .IN1(n30), .IN2(\data_i[1][19] ), .IN3(n14), .IN4(
        \data_i[0][19] ), .Q(n257) );
  AO22X1 U268 ( .IN1(n31), .IN2(\data_i[6][19] ), .IN3(n15), .IN4(
        \data_i[7][19] ), .Q(n256) );
  AO22X1 U269 ( .IN1(n32), .IN2(\data_i[5][19] ), .IN3(n16), .IN4(
        \data_i[4][19] ), .Q(n255) );
  NOR4X0 U270 ( .IN1(n258), .IN2(n257), .IN3(n256), .IN4(n255), .QN(n269) );
  AO22X1 U271 ( .IN1(n17), .IN2(\data_i[26][19] ), .IN3(n1), .IN4(
        \data_i[27][19] ), .Q(n262) );
  AO22X1 U272 ( .IN1(n18), .IN2(\data_i[25][19] ), .IN3(n2), .IN4(
        \data_i[24][19] ), .Q(n261) );
  AO22X1 U273 ( .IN1(n19), .IN2(\data_i[30][19] ), .IN3(n3), .IN4(
        \data_i[31][19] ), .Q(n260) );
  AO22X1 U274 ( .IN1(n20), .IN2(\data_i[29][19] ), .IN3(n4), .IN4(
        \data_i[28][19] ), .Q(n259) );
  NOR4X0 U275 ( .IN1(n262), .IN2(n261), .IN3(n260), .IN4(n259), .QN(n268) );
  AO22X1 U276 ( .IN1(n21), .IN2(\data_i[18][19] ), .IN3(n5), .IN4(
        \data_i[19][19] ), .Q(n266) );
  AO22X1 U277 ( .IN1(n22), .IN2(\data_i[17][19] ), .IN3(n6), .IN4(
        \data_i[16][19] ), .Q(n265) );
  AO22X1 U278 ( .IN1(n23), .IN2(\data_i[22][19] ), .IN3(n7), .IN4(
        \data_i[23][19] ), .Q(n264) );
  AO22X1 U279 ( .IN1(n24), .IN2(\data_i[21][19] ), .IN3(n8), .IN4(
        \data_i[20][19] ), .Q(n263) );
  NOR4X0 U280 ( .IN1(n266), .IN2(n265), .IN3(n264), .IN4(n263), .QN(n267) );
  NAND4X0 U281 ( .IN1(n270), .IN2(n269), .IN3(n268), .IN4(n267), .QN(
        data_o[19]) );
  AO22X1 U282 ( .IN1(n25), .IN2(\data_i[10][1] ), .IN3(n9), .IN4(
        \data_i[11][1] ), .Q(n274) );
  AO22X1 U283 ( .IN1(n26), .IN2(\data_i[9][1] ), .IN3(n10), .IN4(
        \data_i[8][1] ), .Q(n273) );
  AO22X1 U284 ( .IN1(n27), .IN2(\data_i[14][1] ), .IN3(n11), .IN4(
        \data_i[15][1] ), .Q(n272) );
  AO22X1 U285 ( .IN1(n28), .IN2(\data_i[13][1] ), .IN3(n12), .IN4(
        \data_i[12][1] ), .Q(n271) );
  NOR4X0 U286 ( .IN1(n274), .IN2(n273), .IN3(n272), .IN4(n271), .QN(n290) );
  AO22X1 U287 ( .IN1(n29), .IN2(\data_i[2][1] ), .IN3(n13), .IN4(
        \data_i[3][1] ), .Q(n278) );
  AO22X1 U288 ( .IN1(n30), .IN2(\data_i[1][1] ), .IN3(n14), .IN4(
        \data_i[0][1] ), .Q(n277) );
  AO22X1 U289 ( .IN1(n31), .IN2(\data_i[6][1] ), .IN3(n15), .IN4(
        \data_i[7][1] ), .Q(n276) );
  AO22X1 U290 ( .IN1(n32), .IN2(\data_i[5][1] ), .IN3(n16), .IN4(
        \data_i[4][1] ), .Q(n275) );
  NOR4X0 U291 ( .IN1(n278), .IN2(n277), .IN3(n276), .IN4(n275), .QN(n289) );
  AO22X1 U292 ( .IN1(n17), .IN2(\data_i[26][1] ), .IN3(n1), .IN4(
        \data_i[27][1] ), .Q(n282) );
  AO22X1 U293 ( .IN1(n18), .IN2(\data_i[25][1] ), .IN3(n2), .IN4(
        \data_i[24][1] ), .Q(n281) );
  AO22X1 U294 ( .IN1(n19), .IN2(\data_i[30][1] ), .IN3(n3), .IN4(
        \data_i[31][1] ), .Q(n280) );
  AO22X1 U295 ( .IN1(n20), .IN2(\data_i[29][1] ), .IN3(n4), .IN4(
        \data_i[28][1] ), .Q(n279) );
  NOR4X0 U296 ( .IN1(n282), .IN2(n281), .IN3(n280), .IN4(n279), .QN(n288) );
  AO22X1 U297 ( .IN1(n21), .IN2(\data_i[18][1] ), .IN3(n5), .IN4(
        \data_i[19][1] ), .Q(n286) );
  AO22X1 U298 ( .IN1(n22), .IN2(\data_i[17][1] ), .IN3(n6), .IN4(
        \data_i[16][1] ), .Q(n285) );
  AO22X1 U299 ( .IN1(n23), .IN2(\data_i[22][1] ), .IN3(n7), .IN4(
        \data_i[23][1] ), .Q(n284) );
  AO22X1 U300 ( .IN1(n24), .IN2(\data_i[21][1] ), .IN3(n8), .IN4(
        \data_i[20][1] ), .Q(n283) );
  NOR4X0 U301 ( .IN1(n286), .IN2(n285), .IN3(n284), .IN4(n283), .QN(n287) );
  NAND4X0 U302 ( .IN1(n290), .IN2(n289), .IN3(n288), .IN4(n287), .QN(data_o[1]) );
  AO22X1 U303 ( .IN1(n25), .IN2(\data_i[10][20] ), .IN3(n9), .IN4(
        \data_i[11][20] ), .Q(n294) );
  AO22X1 U304 ( .IN1(n26), .IN2(\data_i[9][20] ), .IN3(n10), .IN4(
        \data_i[8][20] ), .Q(n293) );
  AO22X1 U305 ( .IN1(n27), .IN2(\data_i[14][20] ), .IN3(n11), .IN4(
        \data_i[15][20] ), .Q(n292) );
  AO22X1 U306 ( .IN1(n28), .IN2(\data_i[13][20] ), .IN3(n12), .IN4(
        \data_i[12][20] ), .Q(n291) );
  NOR4X0 U307 ( .IN1(n294), .IN2(n293), .IN3(n292), .IN4(n291), .QN(n310) );
  AO22X1 U308 ( .IN1(n29), .IN2(\data_i[2][20] ), .IN3(n13), .IN4(
        \data_i[3][20] ), .Q(n298) );
  AO22X1 U309 ( .IN1(n30), .IN2(\data_i[1][20] ), .IN3(n14), .IN4(
        \data_i[0][20] ), .Q(n297) );
  AO22X1 U310 ( .IN1(n31), .IN2(\data_i[6][20] ), .IN3(n15), .IN4(
        \data_i[7][20] ), .Q(n296) );
  AO22X1 U311 ( .IN1(n32), .IN2(\data_i[5][20] ), .IN3(n16), .IN4(
        \data_i[4][20] ), .Q(n295) );
  NOR4X0 U312 ( .IN1(n298), .IN2(n297), .IN3(n296), .IN4(n295), .QN(n309) );
  AO22X1 U313 ( .IN1(n17), .IN2(\data_i[26][20] ), .IN3(n1), .IN4(
        \data_i[27][20] ), .Q(n302) );
  AO22X1 U314 ( .IN1(n18), .IN2(\data_i[25][20] ), .IN3(n2), .IN4(
        \data_i[24][20] ), .Q(n301) );
  AO22X1 U315 ( .IN1(n19), .IN2(\data_i[30][20] ), .IN3(n3), .IN4(
        \data_i[31][20] ), .Q(n300) );
  AO22X1 U316 ( .IN1(n20), .IN2(\data_i[29][20] ), .IN3(n4), .IN4(
        \data_i[28][20] ), .Q(n299) );
  NOR4X0 U317 ( .IN1(n302), .IN2(n301), .IN3(n300), .IN4(n299), .QN(n308) );
  AO22X1 U318 ( .IN1(n21), .IN2(\data_i[18][20] ), .IN3(n5), .IN4(
        \data_i[19][20] ), .Q(n306) );
  AO22X1 U319 ( .IN1(n22), .IN2(\data_i[17][20] ), .IN3(n6), .IN4(
        \data_i[16][20] ), .Q(n305) );
  AO22X1 U320 ( .IN1(n23), .IN2(\data_i[22][20] ), .IN3(n7), .IN4(
        \data_i[23][20] ), .Q(n304) );
  AO22X1 U321 ( .IN1(n24), .IN2(\data_i[21][20] ), .IN3(n8), .IN4(
        \data_i[20][20] ), .Q(n303) );
  NOR4X0 U322 ( .IN1(n306), .IN2(n305), .IN3(n304), .IN4(n303), .QN(n307) );
  NAND4X0 U323 ( .IN1(n310), .IN2(n309), .IN3(n308), .IN4(n307), .QN(
        data_o[20]) );
  AO22X1 U324 ( .IN1(n25), .IN2(\data_i[10][21] ), .IN3(n9), .IN4(
        \data_i[11][21] ), .Q(n314) );
  AO22X1 U325 ( .IN1(n26), .IN2(\data_i[9][21] ), .IN3(n10), .IN4(
        \data_i[8][21] ), .Q(n313) );
  AO22X1 U326 ( .IN1(n27), .IN2(\data_i[14][21] ), .IN3(n11), .IN4(
        \data_i[15][21] ), .Q(n312) );
  AO22X1 U327 ( .IN1(n28), .IN2(\data_i[13][21] ), .IN3(n12), .IN4(
        \data_i[12][21] ), .Q(n311) );
  NOR4X0 U328 ( .IN1(n314), .IN2(n313), .IN3(n312), .IN4(n311), .QN(n330) );
  AO22X1 U329 ( .IN1(n29), .IN2(\data_i[2][21] ), .IN3(n13), .IN4(
        \data_i[3][21] ), .Q(n318) );
  AO22X1 U330 ( .IN1(n30), .IN2(\data_i[1][21] ), .IN3(n14), .IN4(
        \data_i[0][21] ), .Q(n317) );
  AO22X1 U331 ( .IN1(n31), .IN2(\data_i[6][21] ), .IN3(n15), .IN4(
        \data_i[7][21] ), .Q(n316) );
  AO22X1 U332 ( .IN1(n32), .IN2(\data_i[5][21] ), .IN3(n16), .IN4(
        \data_i[4][21] ), .Q(n315) );
  NOR4X0 U333 ( .IN1(n318), .IN2(n317), .IN3(n316), .IN4(n315), .QN(n329) );
  AO22X1 U334 ( .IN1(n17), .IN2(\data_i[26][21] ), .IN3(n1), .IN4(
        \data_i[27][21] ), .Q(n322) );
  AO22X1 U335 ( .IN1(n18), .IN2(\data_i[25][21] ), .IN3(n2), .IN4(
        \data_i[24][21] ), .Q(n321) );
  AO22X1 U336 ( .IN1(n19), .IN2(\data_i[30][21] ), .IN3(n3), .IN4(
        \data_i[31][21] ), .Q(n320) );
  AO22X1 U337 ( .IN1(n20), .IN2(\data_i[29][21] ), .IN3(n4), .IN4(
        \data_i[28][21] ), .Q(n319) );
  NOR4X0 U338 ( .IN1(n322), .IN2(n321), .IN3(n320), .IN4(n319), .QN(n328) );
  AO22X1 U339 ( .IN1(n21), .IN2(\data_i[18][21] ), .IN3(n5), .IN4(
        \data_i[19][21] ), .Q(n326) );
  AO22X1 U340 ( .IN1(n22), .IN2(\data_i[17][21] ), .IN3(n6), .IN4(
        \data_i[16][21] ), .Q(n325) );
  AO22X1 U341 ( .IN1(n23), .IN2(\data_i[22][21] ), .IN3(n7), .IN4(
        \data_i[23][21] ), .Q(n324) );
  AO22X1 U342 ( .IN1(n24), .IN2(\data_i[21][21] ), .IN3(n8), .IN4(
        \data_i[20][21] ), .Q(n323) );
  NOR4X0 U343 ( .IN1(n326), .IN2(n325), .IN3(n324), .IN4(n323), .QN(n327) );
  NAND4X0 U344 ( .IN1(n330), .IN2(n329), .IN3(n328), .IN4(n327), .QN(
        data_o[21]) );
  AO22X1 U345 ( .IN1(n25), .IN2(\data_i[10][22] ), .IN3(n9), .IN4(
        \data_i[11][22] ), .Q(n334) );
  AO22X1 U346 ( .IN1(n26), .IN2(\data_i[9][22] ), .IN3(n10), .IN4(
        \data_i[8][22] ), .Q(n333) );
  AO22X1 U347 ( .IN1(n27), .IN2(\data_i[14][22] ), .IN3(n11), .IN4(
        \data_i[15][22] ), .Q(n332) );
  AO22X1 U348 ( .IN1(n28), .IN2(\data_i[13][22] ), .IN3(n12), .IN4(
        \data_i[12][22] ), .Q(n331) );
  NOR4X0 U349 ( .IN1(n334), .IN2(n333), .IN3(n332), .IN4(n331), .QN(n350) );
  AO22X1 U350 ( .IN1(n29), .IN2(\data_i[2][22] ), .IN3(n13), .IN4(
        \data_i[3][22] ), .Q(n338) );
  AO22X1 U351 ( .IN1(n30), .IN2(\data_i[1][22] ), .IN3(n14), .IN4(
        \data_i[0][22] ), .Q(n337) );
  AO22X1 U352 ( .IN1(n31), .IN2(\data_i[6][22] ), .IN3(n15), .IN4(
        \data_i[7][22] ), .Q(n336) );
  AO22X1 U353 ( .IN1(n32), .IN2(\data_i[5][22] ), .IN3(n16), .IN4(
        \data_i[4][22] ), .Q(n335) );
  NOR4X0 U354 ( .IN1(n338), .IN2(n337), .IN3(n336), .IN4(n335), .QN(n349) );
  AO22X1 U355 ( .IN1(n17), .IN2(\data_i[26][22] ), .IN3(n1), .IN4(
        \data_i[27][22] ), .Q(n342) );
  AO22X1 U356 ( .IN1(n18), .IN2(\data_i[25][22] ), .IN3(n2), .IN4(
        \data_i[24][22] ), .Q(n341) );
  AO22X1 U357 ( .IN1(n19), .IN2(\data_i[30][22] ), .IN3(n3), .IN4(
        \data_i[31][22] ), .Q(n340) );
  AO22X1 U358 ( .IN1(n20), .IN2(\data_i[29][22] ), .IN3(n4), .IN4(
        \data_i[28][22] ), .Q(n339) );
  NOR4X0 U359 ( .IN1(n342), .IN2(n341), .IN3(n340), .IN4(n339), .QN(n348) );
  AO22X1 U360 ( .IN1(n21), .IN2(\data_i[18][22] ), .IN3(n5), .IN4(
        \data_i[19][22] ), .Q(n346) );
  AO22X1 U361 ( .IN1(n22), .IN2(\data_i[17][22] ), .IN3(n6), .IN4(
        \data_i[16][22] ), .Q(n345) );
  AO22X1 U362 ( .IN1(n23), .IN2(\data_i[22][22] ), .IN3(n7), .IN4(
        \data_i[23][22] ), .Q(n344) );
  AO22X1 U363 ( .IN1(n24), .IN2(\data_i[21][22] ), .IN3(n8), .IN4(
        \data_i[20][22] ), .Q(n343) );
  NOR4X0 U364 ( .IN1(n346), .IN2(n345), .IN3(n344), .IN4(n343), .QN(n347) );
  NAND4X0 U365 ( .IN1(n350), .IN2(n349), .IN3(n348), .IN4(n347), .QN(
        data_o[22]) );
  AO22X1 U366 ( .IN1(n25), .IN2(\data_i[10][23] ), .IN3(n9), .IN4(
        \data_i[11][23] ), .Q(n354) );
  AO22X1 U367 ( .IN1(n26), .IN2(\data_i[9][23] ), .IN3(n10), .IN4(
        \data_i[8][23] ), .Q(n353) );
  AO22X1 U368 ( .IN1(n27), .IN2(\data_i[14][23] ), .IN3(n11), .IN4(
        \data_i[15][23] ), .Q(n352) );
  AO22X1 U369 ( .IN1(n28), .IN2(\data_i[13][23] ), .IN3(n12), .IN4(
        \data_i[12][23] ), .Q(n351) );
  NOR4X0 U370 ( .IN1(n354), .IN2(n353), .IN3(n352), .IN4(n351), .QN(n370) );
  AO22X1 U371 ( .IN1(n29), .IN2(\data_i[2][23] ), .IN3(n13), .IN4(
        \data_i[3][23] ), .Q(n358) );
  AO22X1 U372 ( .IN1(n30), .IN2(\data_i[1][23] ), .IN3(n14), .IN4(
        \data_i[0][23] ), .Q(n357) );
  AO22X1 U373 ( .IN1(n31), .IN2(\data_i[6][23] ), .IN3(n15), .IN4(
        \data_i[7][23] ), .Q(n356) );
  AO22X1 U374 ( .IN1(n32), .IN2(\data_i[5][23] ), .IN3(n16), .IN4(
        \data_i[4][23] ), .Q(n355) );
  NOR4X0 U375 ( .IN1(n358), .IN2(n357), .IN3(n356), .IN4(n355), .QN(n369) );
  AO22X1 U376 ( .IN1(n17), .IN2(\data_i[26][23] ), .IN3(n1), .IN4(
        \data_i[27][23] ), .Q(n362) );
  AO22X1 U377 ( .IN1(n18), .IN2(\data_i[25][23] ), .IN3(n2), .IN4(
        \data_i[24][23] ), .Q(n361) );
  AO22X1 U378 ( .IN1(n19), .IN2(\data_i[30][23] ), .IN3(n3), .IN4(
        \data_i[31][23] ), .Q(n360) );
  AO22X1 U379 ( .IN1(n20), .IN2(\data_i[29][23] ), .IN3(n4), .IN4(
        \data_i[28][23] ), .Q(n359) );
  NOR4X0 U380 ( .IN1(n362), .IN2(n361), .IN3(n360), .IN4(n359), .QN(n368) );
  AO22X1 U381 ( .IN1(n21), .IN2(\data_i[18][23] ), .IN3(n5), .IN4(
        \data_i[19][23] ), .Q(n366) );
  AO22X1 U382 ( .IN1(n22), .IN2(\data_i[17][23] ), .IN3(n6), .IN4(
        \data_i[16][23] ), .Q(n365) );
  AO22X1 U383 ( .IN1(n23), .IN2(\data_i[22][23] ), .IN3(n7), .IN4(
        \data_i[23][23] ), .Q(n364) );
  AO22X1 U384 ( .IN1(n24), .IN2(\data_i[21][23] ), .IN3(n8), .IN4(
        \data_i[20][23] ), .Q(n363) );
  NOR4X0 U385 ( .IN1(n366), .IN2(n365), .IN3(n364), .IN4(n363), .QN(n367) );
  NAND4X0 U386 ( .IN1(n370), .IN2(n369), .IN3(n368), .IN4(n367), .QN(
        data_o[23]) );
  AO22X1 U387 ( .IN1(n25), .IN2(\data_i[10][24] ), .IN3(n9), .IN4(
        \data_i[11][24] ), .Q(n374) );
  AO22X1 U388 ( .IN1(n26), .IN2(\data_i[9][24] ), .IN3(n10), .IN4(
        \data_i[8][24] ), .Q(n373) );
  AO22X1 U389 ( .IN1(n27), .IN2(\data_i[14][24] ), .IN3(n11), .IN4(
        \data_i[15][24] ), .Q(n372) );
  AO22X1 U390 ( .IN1(n28), .IN2(\data_i[13][24] ), .IN3(n12), .IN4(
        \data_i[12][24] ), .Q(n371) );
  NOR4X0 U391 ( .IN1(n374), .IN2(n373), .IN3(n372), .IN4(n371), .QN(n390) );
  AO22X1 U392 ( .IN1(n29), .IN2(\data_i[2][24] ), .IN3(n13), .IN4(
        \data_i[3][24] ), .Q(n378) );
  AO22X1 U393 ( .IN1(n30), .IN2(\data_i[1][24] ), .IN3(n14), .IN4(
        \data_i[0][24] ), .Q(n377) );
  AO22X1 U394 ( .IN1(n31), .IN2(\data_i[6][24] ), .IN3(n15), .IN4(
        \data_i[7][24] ), .Q(n376) );
  AO22X1 U395 ( .IN1(n32), .IN2(\data_i[5][24] ), .IN3(n16), .IN4(
        \data_i[4][24] ), .Q(n375) );
  NOR4X0 U396 ( .IN1(n378), .IN2(n377), .IN3(n376), .IN4(n375), .QN(n389) );
  AO22X1 U397 ( .IN1(n17), .IN2(\data_i[26][24] ), .IN3(n1), .IN4(
        \data_i[27][24] ), .Q(n382) );
  AO22X1 U398 ( .IN1(n18), .IN2(\data_i[25][24] ), .IN3(n2), .IN4(
        \data_i[24][24] ), .Q(n381) );
  AO22X1 U399 ( .IN1(n19), .IN2(\data_i[30][24] ), .IN3(n3), .IN4(
        \data_i[31][24] ), .Q(n380) );
  AO22X1 U400 ( .IN1(n20), .IN2(\data_i[29][24] ), .IN3(n4), .IN4(
        \data_i[28][24] ), .Q(n379) );
  NOR4X0 U401 ( .IN1(n382), .IN2(n381), .IN3(n380), .IN4(n379), .QN(n388) );
  AO22X1 U402 ( .IN1(n21), .IN2(\data_i[18][24] ), .IN3(n5), .IN4(
        \data_i[19][24] ), .Q(n386) );
  AO22X1 U403 ( .IN1(n22), .IN2(\data_i[17][24] ), .IN3(n6), .IN4(
        \data_i[16][24] ), .Q(n385) );
  AO22X1 U404 ( .IN1(n23), .IN2(\data_i[22][24] ), .IN3(n7), .IN4(
        \data_i[23][24] ), .Q(n384) );
  AO22X1 U405 ( .IN1(n24), .IN2(\data_i[21][24] ), .IN3(n8), .IN4(
        \data_i[20][24] ), .Q(n383) );
  NOR4X0 U406 ( .IN1(n386), .IN2(n385), .IN3(n384), .IN4(n383), .QN(n387) );
  NAND4X0 U407 ( .IN1(n390), .IN2(n389), .IN3(n388), .IN4(n387), .QN(
        data_o[24]) );
  AO22X1 U408 ( .IN1(n25), .IN2(\data_i[10][25] ), .IN3(n9), .IN4(
        \data_i[11][25] ), .Q(n394) );
  AO22X1 U409 ( .IN1(n26), .IN2(\data_i[9][25] ), .IN3(n10), .IN4(
        \data_i[8][25] ), .Q(n393) );
  AO22X1 U410 ( .IN1(n27), .IN2(\data_i[14][25] ), .IN3(n11), .IN4(
        \data_i[15][25] ), .Q(n392) );
  AO22X1 U411 ( .IN1(n28), .IN2(\data_i[13][25] ), .IN3(n12), .IN4(
        \data_i[12][25] ), .Q(n391) );
  NOR4X0 U412 ( .IN1(n394), .IN2(n393), .IN3(n392), .IN4(n391), .QN(n410) );
  AO22X1 U413 ( .IN1(n29), .IN2(\data_i[2][25] ), .IN3(n13), .IN4(
        \data_i[3][25] ), .Q(n398) );
  AO22X1 U414 ( .IN1(n30), .IN2(\data_i[1][25] ), .IN3(n14), .IN4(
        \data_i[0][25] ), .Q(n397) );
  AO22X1 U415 ( .IN1(n31), .IN2(\data_i[6][25] ), .IN3(n15), .IN4(
        \data_i[7][25] ), .Q(n396) );
  AO22X1 U416 ( .IN1(n32), .IN2(\data_i[5][25] ), .IN3(n16), .IN4(
        \data_i[4][25] ), .Q(n395) );
  NOR4X0 U417 ( .IN1(n398), .IN2(n397), .IN3(n396), .IN4(n395), .QN(n409) );
  AO22X1 U418 ( .IN1(n17), .IN2(\data_i[26][25] ), .IN3(n1), .IN4(
        \data_i[27][25] ), .Q(n402) );
  AO22X1 U419 ( .IN1(n18), .IN2(\data_i[25][25] ), .IN3(n2), .IN4(
        \data_i[24][25] ), .Q(n401) );
  AO22X1 U420 ( .IN1(n19), .IN2(\data_i[30][25] ), .IN3(n3), .IN4(
        \data_i[31][25] ), .Q(n400) );
  AO22X1 U421 ( .IN1(n20), .IN2(\data_i[29][25] ), .IN3(n4), .IN4(
        \data_i[28][25] ), .Q(n399) );
  NOR4X0 U422 ( .IN1(n402), .IN2(n401), .IN3(n400), .IN4(n399), .QN(n408) );
  AO22X1 U423 ( .IN1(n21), .IN2(\data_i[18][25] ), .IN3(n5), .IN4(
        \data_i[19][25] ), .Q(n406) );
  AO22X1 U424 ( .IN1(n22), .IN2(\data_i[17][25] ), .IN3(n6), .IN4(
        \data_i[16][25] ), .Q(n405) );
  AO22X1 U425 ( .IN1(n23), .IN2(\data_i[22][25] ), .IN3(n7), .IN4(
        \data_i[23][25] ), .Q(n404) );
  AO22X1 U426 ( .IN1(n24), .IN2(\data_i[21][25] ), .IN3(n8), .IN4(
        \data_i[20][25] ), .Q(n403) );
  NOR4X0 U427 ( .IN1(n406), .IN2(n405), .IN3(n404), .IN4(n403), .QN(n407) );
  NAND4X0 U428 ( .IN1(n410), .IN2(n409), .IN3(n408), .IN4(n407), .QN(
        data_o[25]) );
  AO22X1 U429 ( .IN1(n25), .IN2(\data_i[10][26] ), .IN3(n9), .IN4(
        \data_i[11][26] ), .Q(n414) );
  AO22X1 U430 ( .IN1(n26), .IN2(\data_i[9][26] ), .IN3(n10), .IN4(
        \data_i[8][26] ), .Q(n413) );
  AO22X1 U431 ( .IN1(n27), .IN2(\data_i[14][26] ), .IN3(n11), .IN4(
        \data_i[15][26] ), .Q(n412) );
  AO22X1 U432 ( .IN1(n28), .IN2(\data_i[13][26] ), .IN3(n12), .IN4(
        \data_i[12][26] ), .Q(n411) );
  NOR4X0 U433 ( .IN1(n414), .IN2(n413), .IN3(n412), .IN4(n411), .QN(n430) );
  AO22X1 U434 ( .IN1(n29), .IN2(\data_i[2][26] ), .IN3(n13), .IN4(
        \data_i[3][26] ), .Q(n418) );
  AO22X1 U435 ( .IN1(n30), .IN2(\data_i[1][26] ), .IN3(n14), .IN4(
        \data_i[0][26] ), .Q(n417) );
  AO22X1 U436 ( .IN1(n31), .IN2(\data_i[6][26] ), .IN3(n15), .IN4(
        \data_i[7][26] ), .Q(n416) );
  AO22X1 U437 ( .IN1(n32), .IN2(\data_i[5][26] ), .IN3(n16), .IN4(
        \data_i[4][26] ), .Q(n415) );
  NOR4X0 U438 ( .IN1(n418), .IN2(n417), .IN3(n416), .IN4(n415), .QN(n429) );
  AO22X1 U439 ( .IN1(n17), .IN2(\data_i[26][26] ), .IN3(n1), .IN4(
        \data_i[27][26] ), .Q(n422) );
  AO22X1 U440 ( .IN1(n18), .IN2(\data_i[25][26] ), .IN3(n2), .IN4(
        \data_i[24][26] ), .Q(n421) );
  AO22X1 U441 ( .IN1(n19), .IN2(\data_i[30][26] ), .IN3(n3), .IN4(
        \data_i[31][26] ), .Q(n420) );
  AO22X1 U442 ( .IN1(n20), .IN2(\data_i[29][26] ), .IN3(n4), .IN4(
        \data_i[28][26] ), .Q(n419) );
  NOR4X0 U443 ( .IN1(n422), .IN2(n421), .IN3(n420), .IN4(n419), .QN(n428) );
  AO22X1 U444 ( .IN1(n21), .IN2(\data_i[18][26] ), .IN3(n5), .IN4(
        \data_i[19][26] ), .Q(n426) );
  AO22X1 U445 ( .IN1(n22), .IN2(\data_i[17][26] ), .IN3(n6), .IN4(
        \data_i[16][26] ), .Q(n425) );
  AO22X1 U446 ( .IN1(n23), .IN2(\data_i[22][26] ), .IN3(n7), .IN4(
        \data_i[23][26] ), .Q(n424) );
  AO22X1 U447 ( .IN1(n24), .IN2(\data_i[21][26] ), .IN3(n8), .IN4(
        \data_i[20][26] ), .Q(n423) );
  NOR4X0 U448 ( .IN1(n426), .IN2(n425), .IN3(n424), .IN4(n423), .QN(n427) );
  NAND4X0 U449 ( .IN1(n430), .IN2(n429), .IN3(n428), .IN4(n427), .QN(
        data_o[26]) );
  AO22X1 U450 ( .IN1(n25), .IN2(\data_i[10][27] ), .IN3(n9), .IN4(
        \data_i[11][27] ), .Q(n434) );
  AO22X1 U451 ( .IN1(n26), .IN2(\data_i[9][27] ), .IN3(n10), .IN4(
        \data_i[8][27] ), .Q(n433) );
  AO22X1 U452 ( .IN1(n27), .IN2(\data_i[14][27] ), .IN3(n11), .IN4(
        \data_i[15][27] ), .Q(n432) );
  AO22X1 U453 ( .IN1(n28), .IN2(\data_i[13][27] ), .IN3(n12), .IN4(
        \data_i[12][27] ), .Q(n431) );
  NOR4X0 U454 ( .IN1(n434), .IN2(n433), .IN3(n432), .IN4(n431), .QN(n450) );
  AO22X1 U455 ( .IN1(n29), .IN2(\data_i[2][27] ), .IN3(n13), .IN4(
        \data_i[3][27] ), .Q(n438) );
  AO22X1 U456 ( .IN1(n30), .IN2(\data_i[1][27] ), .IN3(n14), .IN4(
        \data_i[0][27] ), .Q(n437) );
  AO22X1 U457 ( .IN1(n31), .IN2(\data_i[6][27] ), .IN3(n15), .IN4(
        \data_i[7][27] ), .Q(n436) );
  AO22X1 U458 ( .IN1(n32), .IN2(\data_i[5][27] ), .IN3(n16), .IN4(
        \data_i[4][27] ), .Q(n435) );
  NOR4X0 U459 ( .IN1(n438), .IN2(n437), .IN3(n436), .IN4(n435), .QN(n449) );
  AO22X1 U460 ( .IN1(n17), .IN2(\data_i[26][27] ), .IN3(n1), .IN4(
        \data_i[27][27] ), .Q(n442) );
  AO22X1 U461 ( .IN1(n18), .IN2(\data_i[25][27] ), .IN3(n2), .IN4(
        \data_i[24][27] ), .Q(n441) );
  AO22X1 U462 ( .IN1(n19), .IN2(\data_i[30][27] ), .IN3(n3), .IN4(
        \data_i[31][27] ), .Q(n440) );
  AO22X1 U463 ( .IN1(n20), .IN2(\data_i[29][27] ), .IN3(n4), .IN4(
        \data_i[28][27] ), .Q(n439) );
  NOR4X0 U464 ( .IN1(n442), .IN2(n441), .IN3(n440), .IN4(n439), .QN(n448) );
  AO22X1 U465 ( .IN1(n21), .IN2(\data_i[18][27] ), .IN3(n5), .IN4(
        \data_i[19][27] ), .Q(n446) );
  AO22X1 U466 ( .IN1(n22), .IN2(\data_i[17][27] ), .IN3(n6), .IN4(
        \data_i[16][27] ), .Q(n445) );
  AO22X1 U467 ( .IN1(n23), .IN2(\data_i[22][27] ), .IN3(n7), .IN4(
        \data_i[23][27] ), .Q(n444) );
  AO22X1 U468 ( .IN1(n24), .IN2(\data_i[21][27] ), .IN3(n8), .IN4(
        \data_i[20][27] ), .Q(n443) );
  NOR4X0 U469 ( .IN1(n446), .IN2(n445), .IN3(n444), .IN4(n443), .QN(n447) );
  NAND4X0 U470 ( .IN1(n450), .IN2(n449), .IN3(n448), .IN4(n447), .QN(
        data_o[27]) );
  AO22X1 U471 ( .IN1(n25), .IN2(\data_i[10][28] ), .IN3(n9), .IN4(
        \data_i[11][28] ), .Q(n454) );
  AO22X1 U472 ( .IN1(n26), .IN2(\data_i[9][28] ), .IN3(n10), .IN4(
        \data_i[8][28] ), .Q(n453) );
  AO22X1 U473 ( .IN1(n27), .IN2(\data_i[14][28] ), .IN3(n11), .IN4(
        \data_i[15][28] ), .Q(n452) );
  AO22X1 U474 ( .IN1(n28), .IN2(\data_i[13][28] ), .IN3(n12), .IN4(
        \data_i[12][28] ), .Q(n451) );
  NOR4X0 U475 ( .IN1(n454), .IN2(n453), .IN3(n452), .IN4(n451), .QN(n470) );
  AO22X1 U476 ( .IN1(n29), .IN2(\data_i[2][28] ), .IN3(n13), .IN4(
        \data_i[3][28] ), .Q(n458) );
  AO22X1 U477 ( .IN1(n30), .IN2(\data_i[1][28] ), .IN3(n14), .IN4(
        \data_i[0][28] ), .Q(n457) );
  AO22X1 U478 ( .IN1(n31), .IN2(\data_i[6][28] ), .IN3(n15), .IN4(
        \data_i[7][28] ), .Q(n456) );
  AO22X1 U479 ( .IN1(n32), .IN2(\data_i[5][28] ), .IN3(n16), .IN4(
        \data_i[4][28] ), .Q(n455) );
  NOR4X0 U480 ( .IN1(n458), .IN2(n457), .IN3(n456), .IN4(n455), .QN(n469) );
  AO22X1 U481 ( .IN1(n17), .IN2(\data_i[26][28] ), .IN3(n1), .IN4(
        \data_i[27][28] ), .Q(n462) );
  AO22X1 U482 ( .IN1(n18), .IN2(\data_i[25][28] ), .IN3(n2), .IN4(
        \data_i[24][28] ), .Q(n461) );
  AO22X1 U483 ( .IN1(n19), .IN2(\data_i[30][28] ), .IN3(n3), .IN4(
        \data_i[31][28] ), .Q(n460) );
  AO22X1 U484 ( .IN1(n20), .IN2(\data_i[29][28] ), .IN3(n4), .IN4(
        \data_i[28][28] ), .Q(n459) );
  NOR4X0 U485 ( .IN1(n462), .IN2(n461), .IN3(n460), .IN4(n459), .QN(n468) );
  AO22X1 U486 ( .IN1(n21), .IN2(\data_i[18][28] ), .IN3(n5), .IN4(
        \data_i[19][28] ), .Q(n466) );
  AO22X1 U487 ( .IN1(n22), .IN2(\data_i[17][28] ), .IN3(n6), .IN4(
        \data_i[16][28] ), .Q(n465) );
  AO22X1 U488 ( .IN1(n23), .IN2(\data_i[22][28] ), .IN3(n7), .IN4(
        \data_i[23][28] ), .Q(n464) );
  AO22X1 U489 ( .IN1(n24), .IN2(\data_i[21][28] ), .IN3(n8), .IN4(
        \data_i[20][28] ), .Q(n463) );
  NOR4X0 U490 ( .IN1(n466), .IN2(n465), .IN3(n464), .IN4(n463), .QN(n467) );
  NAND4X0 U491 ( .IN1(n470), .IN2(n469), .IN3(n468), .IN4(n467), .QN(
        data_o[28]) );
  AO22X1 U492 ( .IN1(n25), .IN2(\data_i[10][29] ), .IN3(n9), .IN4(
        \data_i[11][29] ), .Q(n474) );
  AO22X1 U493 ( .IN1(n26), .IN2(\data_i[9][29] ), .IN3(n10), .IN4(
        \data_i[8][29] ), .Q(n473) );
  AO22X1 U494 ( .IN1(n27), .IN2(\data_i[14][29] ), .IN3(n11), .IN4(
        \data_i[15][29] ), .Q(n472) );
  AO22X1 U495 ( .IN1(n28), .IN2(\data_i[13][29] ), .IN3(n12), .IN4(
        \data_i[12][29] ), .Q(n471) );
  NOR4X0 U496 ( .IN1(n474), .IN2(n473), .IN3(n472), .IN4(n471), .QN(n490) );
  AO22X1 U497 ( .IN1(n29), .IN2(\data_i[2][29] ), .IN3(n13), .IN4(
        \data_i[3][29] ), .Q(n478) );
  AO22X1 U498 ( .IN1(n30), .IN2(\data_i[1][29] ), .IN3(n14), .IN4(
        \data_i[0][29] ), .Q(n477) );
  AO22X1 U499 ( .IN1(n31), .IN2(\data_i[6][29] ), .IN3(n15), .IN4(
        \data_i[7][29] ), .Q(n476) );
  AO22X1 U500 ( .IN1(n32), .IN2(\data_i[5][29] ), .IN3(n16), .IN4(
        \data_i[4][29] ), .Q(n475) );
  NOR4X0 U501 ( .IN1(n478), .IN2(n477), .IN3(n476), .IN4(n475), .QN(n489) );
  AO22X1 U502 ( .IN1(n17), .IN2(\data_i[26][29] ), .IN3(n1), .IN4(
        \data_i[27][29] ), .Q(n482) );
  AO22X1 U503 ( .IN1(n18), .IN2(\data_i[25][29] ), .IN3(n2), .IN4(
        \data_i[24][29] ), .Q(n481) );
  AO22X1 U504 ( .IN1(n19), .IN2(\data_i[30][29] ), .IN3(n3), .IN4(
        \data_i[31][29] ), .Q(n480) );
  AO22X1 U505 ( .IN1(n20), .IN2(\data_i[29][29] ), .IN3(n4), .IN4(
        \data_i[28][29] ), .Q(n479) );
  NOR4X0 U506 ( .IN1(n482), .IN2(n481), .IN3(n480), .IN4(n479), .QN(n488) );
  AO22X1 U507 ( .IN1(n21), .IN2(\data_i[18][29] ), .IN3(n5), .IN4(
        \data_i[19][29] ), .Q(n486) );
  AO22X1 U508 ( .IN1(n22), .IN2(\data_i[17][29] ), .IN3(n6), .IN4(
        \data_i[16][29] ), .Q(n485) );
  AO22X1 U509 ( .IN1(n23), .IN2(\data_i[22][29] ), .IN3(n7), .IN4(
        \data_i[23][29] ), .Q(n484) );
  AO22X1 U510 ( .IN1(n24), .IN2(\data_i[21][29] ), .IN3(n8), .IN4(
        \data_i[20][29] ), .Q(n483) );
  NOR4X0 U511 ( .IN1(n486), .IN2(n485), .IN3(n484), .IN4(n483), .QN(n487) );
  NAND4X0 U512 ( .IN1(n490), .IN2(n489), .IN3(n488), .IN4(n487), .QN(
        data_o[29]) );
  AO22X1 U513 ( .IN1(n25), .IN2(\data_i[10][2] ), .IN3(n9), .IN4(
        \data_i[11][2] ), .Q(n494) );
  AO22X1 U514 ( .IN1(n26), .IN2(\data_i[9][2] ), .IN3(n10), .IN4(
        \data_i[8][2] ), .Q(n493) );
  AO22X1 U515 ( .IN1(n27), .IN2(\data_i[14][2] ), .IN3(n11), .IN4(
        \data_i[15][2] ), .Q(n492) );
  AO22X1 U516 ( .IN1(n28), .IN2(\data_i[13][2] ), .IN3(n12), .IN4(
        \data_i[12][2] ), .Q(n491) );
  NOR4X0 U517 ( .IN1(n494), .IN2(n493), .IN3(n492), .IN4(n491), .QN(n510) );
  AO22X1 U518 ( .IN1(n29), .IN2(\data_i[2][2] ), .IN3(n13), .IN4(
        \data_i[3][2] ), .Q(n498) );
  AO22X1 U519 ( .IN1(n30), .IN2(\data_i[1][2] ), .IN3(n14), .IN4(
        \data_i[0][2] ), .Q(n497) );
  AO22X1 U520 ( .IN1(n31), .IN2(\data_i[6][2] ), .IN3(n15), .IN4(
        \data_i[7][2] ), .Q(n496) );
  AO22X1 U521 ( .IN1(n32), .IN2(\data_i[5][2] ), .IN3(n16), .IN4(
        \data_i[4][2] ), .Q(n495) );
  NOR4X0 U522 ( .IN1(n498), .IN2(n497), .IN3(n496), .IN4(n495), .QN(n509) );
  AO22X1 U523 ( .IN1(n17), .IN2(\data_i[26][2] ), .IN3(n1), .IN4(
        \data_i[27][2] ), .Q(n502) );
  AO22X1 U524 ( .IN1(n18), .IN2(\data_i[25][2] ), .IN3(n2), .IN4(
        \data_i[24][2] ), .Q(n501) );
  AO22X1 U525 ( .IN1(n19), .IN2(\data_i[30][2] ), .IN3(n3), .IN4(
        \data_i[31][2] ), .Q(n500) );
  AO22X1 U526 ( .IN1(n20), .IN2(\data_i[29][2] ), .IN3(n4), .IN4(
        \data_i[28][2] ), .Q(n499) );
  NOR4X0 U527 ( .IN1(n502), .IN2(n501), .IN3(n500), .IN4(n499), .QN(n508) );
  AO22X1 U528 ( .IN1(n21), .IN2(\data_i[18][2] ), .IN3(n5), .IN4(
        \data_i[19][2] ), .Q(n506) );
  AO22X1 U529 ( .IN1(n22), .IN2(\data_i[17][2] ), .IN3(n6), .IN4(
        \data_i[16][2] ), .Q(n505) );
  AO22X1 U530 ( .IN1(n23), .IN2(\data_i[22][2] ), .IN3(n7), .IN4(
        \data_i[23][2] ), .Q(n504) );
  AO22X1 U531 ( .IN1(n24), .IN2(\data_i[21][2] ), .IN3(n8), .IN4(
        \data_i[20][2] ), .Q(n503) );
  NOR4X0 U532 ( .IN1(n506), .IN2(n505), .IN3(n504), .IN4(n503), .QN(n507) );
  NAND4X0 U533 ( .IN1(n510), .IN2(n509), .IN3(n508), .IN4(n507), .QN(data_o[2]) );
  AO22X1 U534 ( .IN1(n25), .IN2(\data_i[10][30] ), .IN3(n9), .IN4(
        \data_i[11][30] ), .Q(n514) );
  AO22X1 U535 ( .IN1(n26), .IN2(\data_i[9][30] ), .IN3(n10), .IN4(
        \data_i[8][30] ), .Q(n513) );
  AO22X1 U536 ( .IN1(n27), .IN2(\data_i[14][30] ), .IN3(n11), .IN4(
        \data_i[15][30] ), .Q(n512) );
  AO22X1 U537 ( .IN1(n28), .IN2(\data_i[13][30] ), .IN3(n12), .IN4(
        \data_i[12][30] ), .Q(n511) );
  NOR4X0 U538 ( .IN1(n514), .IN2(n513), .IN3(n512), .IN4(n511), .QN(n530) );
  AO22X1 U539 ( .IN1(n29), .IN2(\data_i[2][30] ), .IN3(n13), .IN4(
        \data_i[3][30] ), .Q(n518) );
  AO22X1 U540 ( .IN1(n30), .IN2(\data_i[1][30] ), .IN3(n14), .IN4(
        \data_i[0][30] ), .Q(n517) );
  AO22X1 U541 ( .IN1(n31), .IN2(\data_i[6][30] ), .IN3(n15), .IN4(
        \data_i[7][30] ), .Q(n516) );
  AO22X1 U542 ( .IN1(n32), .IN2(\data_i[5][30] ), .IN3(n16), .IN4(
        \data_i[4][30] ), .Q(n515) );
  NOR4X0 U543 ( .IN1(n518), .IN2(n517), .IN3(n516), .IN4(n515), .QN(n529) );
  AO22X1 U544 ( .IN1(n17), .IN2(\data_i[26][30] ), .IN3(n1), .IN4(
        \data_i[27][30] ), .Q(n522) );
  AO22X1 U545 ( .IN1(n18), .IN2(\data_i[25][30] ), .IN3(n2), .IN4(
        \data_i[24][30] ), .Q(n521) );
  AO22X1 U546 ( .IN1(n19), .IN2(\data_i[30][30] ), .IN3(n3), .IN4(
        \data_i[31][30] ), .Q(n520) );
  AO22X1 U547 ( .IN1(n20), .IN2(\data_i[29][30] ), .IN3(n4), .IN4(
        \data_i[28][30] ), .Q(n519) );
  NOR4X0 U548 ( .IN1(n522), .IN2(n521), .IN3(n520), .IN4(n519), .QN(n528) );
  AO22X1 U549 ( .IN1(n21), .IN2(\data_i[18][30] ), .IN3(n5), .IN4(
        \data_i[19][30] ), .Q(n526) );
  AO22X1 U550 ( .IN1(n22), .IN2(\data_i[17][30] ), .IN3(n6), .IN4(
        \data_i[16][30] ), .Q(n525) );
  AO22X1 U551 ( .IN1(n23), .IN2(\data_i[22][30] ), .IN3(n7), .IN4(
        \data_i[23][30] ), .Q(n524) );
  AO22X1 U552 ( .IN1(n24), .IN2(\data_i[21][30] ), .IN3(n8), .IN4(
        \data_i[20][30] ), .Q(n523) );
  NOR4X0 U553 ( .IN1(n526), .IN2(n525), .IN3(n524), .IN4(n523), .QN(n527) );
  NAND4X0 U554 ( .IN1(n530), .IN2(n529), .IN3(n528), .IN4(n527), .QN(
        data_o[30]) );
  AO22X1 U555 ( .IN1(n25), .IN2(\data_i[10][31] ), .IN3(n9), .IN4(
        \data_i[11][31] ), .Q(n534) );
  AO22X1 U556 ( .IN1(n26), .IN2(\data_i[9][31] ), .IN3(n10), .IN4(
        \data_i[8][31] ), .Q(n533) );
  AO22X1 U557 ( .IN1(n27), .IN2(\data_i[14][31] ), .IN3(n11), .IN4(
        \data_i[15][31] ), .Q(n532) );
  AO22X1 U558 ( .IN1(n28), .IN2(\data_i[13][31] ), .IN3(n12), .IN4(
        \data_i[12][31] ), .Q(n531) );
  NOR4X0 U559 ( .IN1(n534), .IN2(n533), .IN3(n532), .IN4(n531), .QN(n550) );
  AO22X1 U560 ( .IN1(n29), .IN2(\data_i[2][31] ), .IN3(n13), .IN4(
        \data_i[3][31] ), .Q(n538) );
  AO22X1 U561 ( .IN1(n30), .IN2(\data_i[1][31] ), .IN3(n14), .IN4(
        \data_i[0][31] ), .Q(n537) );
  AO22X1 U562 ( .IN1(n31), .IN2(\data_i[6][31] ), .IN3(n15), .IN4(
        \data_i[7][31] ), .Q(n536) );
  AO22X1 U563 ( .IN1(n32), .IN2(\data_i[5][31] ), .IN3(n16), .IN4(
        \data_i[4][31] ), .Q(n535) );
  NOR4X0 U564 ( .IN1(n538), .IN2(n537), .IN3(n536), .IN4(n535), .QN(n549) );
  AO22X1 U565 ( .IN1(n17), .IN2(\data_i[26][31] ), .IN3(n1), .IN4(
        \data_i[27][31] ), .Q(n542) );
  AO22X1 U566 ( .IN1(n18), .IN2(\data_i[25][31] ), .IN3(n2), .IN4(
        \data_i[24][31] ), .Q(n541) );
  AO22X1 U567 ( .IN1(n19), .IN2(\data_i[30][31] ), .IN3(n3), .IN4(
        \data_i[31][31] ), .Q(n540) );
  AO22X1 U568 ( .IN1(n20), .IN2(\data_i[29][31] ), .IN3(n4), .IN4(
        \data_i[28][31] ), .Q(n539) );
  NOR4X0 U569 ( .IN1(n542), .IN2(n541), .IN3(n540), .IN4(n539), .QN(n548) );
  AO22X1 U570 ( .IN1(n21), .IN2(\data_i[18][31] ), .IN3(n5), .IN4(
        \data_i[19][31] ), .Q(n546) );
  AO22X1 U571 ( .IN1(n22), .IN2(\data_i[17][31] ), .IN3(n6), .IN4(
        \data_i[16][31] ), .Q(n545) );
  AO22X1 U572 ( .IN1(n23), .IN2(\data_i[22][31] ), .IN3(n7), .IN4(
        \data_i[23][31] ), .Q(n544) );
  AO22X1 U573 ( .IN1(n24), .IN2(\data_i[21][31] ), .IN3(n8), .IN4(
        \data_i[20][31] ), .Q(n543) );
  NOR4X0 U574 ( .IN1(n546), .IN2(n545), .IN3(n544), .IN4(n543), .QN(n547) );
  NAND4X0 U575 ( .IN1(n550), .IN2(n549), .IN3(n548), .IN4(n547), .QN(
        data_o[31]) );
  AO22X1 U576 ( .IN1(n25), .IN2(\data_i[10][3] ), .IN3(n9), .IN4(
        \data_i[11][3] ), .Q(n554) );
  AO22X1 U577 ( .IN1(n26), .IN2(\data_i[9][3] ), .IN3(n10), .IN4(
        \data_i[8][3] ), .Q(n553) );
  AO22X1 U578 ( .IN1(n27), .IN2(\data_i[14][3] ), .IN3(n11), .IN4(
        \data_i[15][3] ), .Q(n552) );
  AO22X1 U579 ( .IN1(n28), .IN2(\data_i[13][3] ), .IN3(n12), .IN4(
        \data_i[12][3] ), .Q(n551) );
  NOR4X0 U580 ( .IN1(n554), .IN2(n553), .IN3(n552), .IN4(n551), .QN(n570) );
  AO22X1 U581 ( .IN1(n29), .IN2(\data_i[2][3] ), .IN3(n13), .IN4(
        \data_i[3][3] ), .Q(n558) );
  AO22X1 U582 ( .IN1(n30), .IN2(\data_i[1][3] ), .IN3(n14), .IN4(
        \data_i[0][3] ), .Q(n557) );
  AO22X1 U583 ( .IN1(n31), .IN2(\data_i[6][3] ), .IN3(n15), .IN4(
        \data_i[7][3] ), .Q(n556) );
  AO22X1 U584 ( .IN1(n32), .IN2(\data_i[5][3] ), .IN3(n16), .IN4(
        \data_i[4][3] ), .Q(n555) );
  NOR4X0 U585 ( .IN1(n558), .IN2(n557), .IN3(n556), .IN4(n555), .QN(n569) );
  AO22X1 U586 ( .IN1(n17), .IN2(\data_i[26][3] ), .IN3(n1), .IN4(
        \data_i[27][3] ), .Q(n562) );
  AO22X1 U587 ( .IN1(n18), .IN2(\data_i[25][3] ), .IN3(n2), .IN4(
        \data_i[24][3] ), .Q(n561) );
  AO22X1 U588 ( .IN1(n19), .IN2(\data_i[30][3] ), .IN3(n3), .IN4(
        \data_i[31][3] ), .Q(n560) );
  AO22X1 U589 ( .IN1(n20), .IN2(\data_i[29][3] ), .IN3(n4), .IN4(
        \data_i[28][3] ), .Q(n559) );
  NOR4X0 U590 ( .IN1(n562), .IN2(n561), .IN3(n560), .IN4(n559), .QN(n568) );
  AO22X1 U591 ( .IN1(n21), .IN2(\data_i[18][3] ), .IN3(n5), .IN4(
        \data_i[19][3] ), .Q(n566) );
  AO22X1 U592 ( .IN1(n22), .IN2(\data_i[17][3] ), .IN3(n6), .IN4(
        \data_i[16][3] ), .Q(n565) );
  AO22X1 U593 ( .IN1(n23), .IN2(\data_i[22][3] ), .IN3(n7), .IN4(
        \data_i[23][3] ), .Q(n564) );
  AO22X1 U594 ( .IN1(n24), .IN2(\data_i[21][3] ), .IN3(n8), .IN4(
        \data_i[20][3] ), .Q(n563) );
  NOR4X0 U595 ( .IN1(n566), .IN2(n565), .IN3(n564), .IN4(n563), .QN(n567) );
  NAND4X0 U596 ( .IN1(n570), .IN2(n569), .IN3(n568), .IN4(n567), .QN(data_o[3]) );
  AO22X1 U597 ( .IN1(n25), .IN2(\data_i[10][4] ), .IN3(n9), .IN4(
        \data_i[11][4] ), .Q(n574) );
  AO22X1 U598 ( .IN1(n26), .IN2(\data_i[9][4] ), .IN3(n10), .IN4(
        \data_i[8][4] ), .Q(n573) );
  AO22X1 U599 ( .IN1(n27), .IN2(\data_i[14][4] ), .IN3(n11), .IN4(
        \data_i[15][4] ), .Q(n572) );
  AO22X1 U600 ( .IN1(n28), .IN2(\data_i[13][4] ), .IN3(n12), .IN4(
        \data_i[12][4] ), .Q(n571) );
  NOR4X0 U601 ( .IN1(n574), .IN2(n573), .IN3(n572), .IN4(n571), .QN(n590) );
  AO22X1 U602 ( .IN1(n29), .IN2(\data_i[2][4] ), .IN3(n13), .IN4(
        \data_i[3][4] ), .Q(n578) );
  AO22X1 U603 ( .IN1(n30), .IN2(\data_i[1][4] ), .IN3(n14), .IN4(
        \data_i[0][4] ), .Q(n577) );
  AO22X1 U604 ( .IN1(n31), .IN2(\data_i[6][4] ), .IN3(n15), .IN4(
        \data_i[7][4] ), .Q(n576) );
  AO22X1 U605 ( .IN1(n32), .IN2(\data_i[5][4] ), .IN3(n16), .IN4(
        \data_i[4][4] ), .Q(n575) );
  NOR4X0 U606 ( .IN1(n578), .IN2(n577), .IN3(n576), .IN4(n575), .QN(n589) );
  AO22X1 U607 ( .IN1(n17), .IN2(\data_i[26][4] ), .IN3(n1), .IN4(
        \data_i[27][4] ), .Q(n582) );
  AO22X1 U608 ( .IN1(n18), .IN2(\data_i[25][4] ), .IN3(n2), .IN4(
        \data_i[24][4] ), .Q(n581) );
  AO22X1 U609 ( .IN1(n19), .IN2(\data_i[30][4] ), .IN3(n3), .IN4(
        \data_i[31][4] ), .Q(n580) );
  AO22X1 U610 ( .IN1(n20), .IN2(\data_i[29][4] ), .IN3(n4), .IN4(
        \data_i[28][4] ), .Q(n579) );
  NOR4X0 U611 ( .IN1(n582), .IN2(n581), .IN3(n580), .IN4(n579), .QN(n588) );
  AO22X1 U612 ( .IN1(n21), .IN2(\data_i[18][4] ), .IN3(n5), .IN4(
        \data_i[19][4] ), .Q(n586) );
  AO22X1 U613 ( .IN1(n22), .IN2(\data_i[17][4] ), .IN3(n6), .IN4(
        \data_i[16][4] ), .Q(n585) );
  AO22X1 U614 ( .IN1(n23), .IN2(\data_i[22][4] ), .IN3(n7), .IN4(
        \data_i[23][4] ), .Q(n584) );
  AO22X1 U615 ( .IN1(n24), .IN2(\data_i[21][4] ), .IN3(n8), .IN4(
        \data_i[20][4] ), .Q(n583) );
  NOR4X0 U616 ( .IN1(n586), .IN2(n585), .IN3(n584), .IN4(n583), .QN(n587) );
  NAND4X0 U617 ( .IN1(n590), .IN2(n589), .IN3(n588), .IN4(n587), .QN(data_o[4]) );
  AO22X1 U618 ( .IN1(n25), .IN2(\data_i[10][5] ), .IN3(n9), .IN4(
        \data_i[11][5] ), .Q(n594) );
  AO22X1 U619 ( .IN1(n26), .IN2(\data_i[9][5] ), .IN3(n10), .IN4(
        \data_i[8][5] ), .Q(n593) );
  AO22X1 U620 ( .IN1(n27), .IN2(\data_i[14][5] ), .IN3(n11), .IN4(
        \data_i[15][5] ), .Q(n592) );
  AO22X1 U621 ( .IN1(n28), .IN2(\data_i[13][5] ), .IN3(n12), .IN4(
        \data_i[12][5] ), .Q(n591) );
  NOR4X0 U622 ( .IN1(n594), .IN2(n593), .IN3(n592), .IN4(n591), .QN(n610) );
  AO22X1 U623 ( .IN1(n29), .IN2(\data_i[2][5] ), .IN3(n13), .IN4(
        \data_i[3][5] ), .Q(n598) );
  AO22X1 U624 ( .IN1(n30), .IN2(\data_i[1][5] ), .IN3(n14), .IN4(
        \data_i[0][5] ), .Q(n597) );
  AO22X1 U625 ( .IN1(n31), .IN2(\data_i[6][5] ), .IN3(n15), .IN4(
        \data_i[7][5] ), .Q(n596) );
  AO22X1 U626 ( .IN1(n32), .IN2(\data_i[5][5] ), .IN3(n16), .IN4(
        \data_i[4][5] ), .Q(n595) );
  NOR4X0 U627 ( .IN1(n598), .IN2(n597), .IN3(n596), .IN4(n595), .QN(n609) );
  AO22X1 U628 ( .IN1(n17), .IN2(\data_i[26][5] ), .IN3(n1), .IN4(
        \data_i[27][5] ), .Q(n602) );
  AO22X1 U629 ( .IN1(n18), .IN2(\data_i[25][5] ), .IN3(n2), .IN4(
        \data_i[24][5] ), .Q(n601) );
  AO22X1 U630 ( .IN1(n19), .IN2(\data_i[30][5] ), .IN3(n3), .IN4(
        \data_i[31][5] ), .Q(n600) );
  AO22X1 U631 ( .IN1(n20), .IN2(\data_i[29][5] ), .IN3(n4), .IN4(
        \data_i[28][5] ), .Q(n599) );
  NOR4X0 U632 ( .IN1(n602), .IN2(n601), .IN3(n600), .IN4(n599), .QN(n608) );
  AO22X1 U633 ( .IN1(n21), .IN2(\data_i[18][5] ), .IN3(n5), .IN4(
        \data_i[19][5] ), .Q(n606) );
  AO22X1 U634 ( .IN1(n22), .IN2(\data_i[17][5] ), .IN3(n6), .IN4(
        \data_i[16][5] ), .Q(n605) );
  AO22X1 U635 ( .IN1(n23), .IN2(\data_i[22][5] ), .IN3(n7), .IN4(
        \data_i[23][5] ), .Q(n604) );
  AO22X1 U636 ( .IN1(n24), .IN2(\data_i[21][5] ), .IN3(n8), .IN4(
        \data_i[20][5] ), .Q(n603) );
  NOR4X0 U637 ( .IN1(n606), .IN2(n605), .IN3(n604), .IN4(n603), .QN(n607) );
  NAND4X0 U638 ( .IN1(n610), .IN2(n609), .IN3(n608), .IN4(n607), .QN(data_o[5]) );
  AO22X1 U639 ( .IN1(n25), .IN2(\data_i[10][6] ), .IN3(n9), .IN4(
        \data_i[11][6] ), .Q(n614) );
  AO22X1 U640 ( .IN1(n26), .IN2(\data_i[9][6] ), .IN3(n10), .IN4(
        \data_i[8][6] ), .Q(n613) );
  AO22X1 U641 ( .IN1(n27), .IN2(\data_i[14][6] ), .IN3(n11), .IN4(
        \data_i[15][6] ), .Q(n612) );
  AO22X1 U642 ( .IN1(n28), .IN2(\data_i[13][6] ), .IN3(n12), .IN4(
        \data_i[12][6] ), .Q(n611) );
  NOR4X0 U643 ( .IN1(n614), .IN2(n613), .IN3(n612), .IN4(n611), .QN(n630) );
  AO22X1 U644 ( .IN1(n29), .IN2(\data_i[2][6] ), .IN3(n13), .IN4(
        \data_i[3][6] ), .Q(n618) );
  AO22X1 U645 ( .IN1(n30), .IN2(\data_i[1][6] ), .IN3(n14), .IN4(
        \data_i[0][6] ), .Q(n617) );
  AO22X1 U646 ( .IN1(n31), .IN2(\data_i[6][6] ), .IN3(n15), .IN4(
        \data_i[7][6] ), .Q(n616) );
  AO22X1 U647 ( .IN1(n32), .IN2(\data_i[5][6] ), .IN3(n16), .IN4(
        \data_i[4][6] ), .Q(n615) );
  NOR4X0 U648 ( .IN1(n618), .IN2(n617), .IN3(n616), .IN4(n615), .QN(n629) );
  AO22X1 U649 ( .IN1(n17), .IN2(\data_i[26][6] ), .IN3(n1), .IN4(
        \data_i[27][6] ), .Q(n622) );
  AO22X1 U650 ( .IN1(n18), .IN2(\data_i[25][6] ), .IN3(n2), .IN4(
        \data_i[24][6] ), .Q(n621) );
  AO22X1 U651 ( .IN1(n19), .IN2(\data_i[30][6] ), .IN3(n3), .IN4(
        \data_i[31][6] ), .Q(n620) );
  AO22X1 U652 ( .IN1(n20), .IN2(\data_i[29][6] ), .IN3(n4), .IN4(
        \data_i[28][6] ), .Q(n619) );
  NOR4X0 U653 ( .IN1(n622), .IN2(n621), .IN3(n620), .IN4(n619), .QN(n628) );
  AO22X1 U654 ( .IN1(n21), .IN2(\data_i[18][6] ), .IN3(n5), .IN4(
        \data_i[19][6] ), .Q(n626) );
  AO22X1 U655 ( .IN1(n22), .IN2(\data_i[17][6] ), .IN3(n6), .IN4(
        \data_i[16][6] ), .Q(n625) );
  AO22X1 U656 ( .IN1(n23), .IN2(\data_i[22][6] ), .IN3(n7), .IN4(
        \data_i[23][6] ), .Q(n624) );
  AO22X1 U657 ( .IN1(n24), .IN2(\data_i[21][6] ), .IN3(n8), .IN4(
        \data_i[20][6] ), .Q(n623) );
  NOR4X0 U658 ( .IN1(n626), .IN2(n625), .IN3(n624), .IN4(n623), .QN(n627) );
  NAND4X0 U659 ( .IN1(n630), .IN2(n629), .IN3(n628), .IN4(n627), .QN(data_o[6]) );
  AO22X1 U660 ( .IN1(n25), .IN2(\data_i[10][7] ), .IN3(n9), .IN4(
        \data_i[11][7] ), .Q(n634) );
  AO22X1 U661 ( .IN1(n26), .IN2(\data_i[9][7] ), .IN3(n10), .IN4(
        \data_i[8][7] ), .Q(n633) );
  AO22X1 U662 ( .IN1(n27), .IN2(\data_i[14][7] ), .IN3(n11), .IN4(
        \data_i[15][7] ), .Q(n632) );
  AO22X1 U663 ( .IN1(n28), .IN2(\data_i[13][7] ), .IN3(n12), .IN4(
        \data_i[12][7] ), .Q(n631) );
  NOR4X0 U664 ( .IN1(n634), .IN2(n633), .IN3(n632), .IN4(n631), .QN(n650) );
  AO22X1 U665 ( .IN1(n29), .IN2(\data_i[2][7] ), .IN3(n13), .IN4(
        \data_i[3][7] ), .Q(n638) );
  AO22X1 U666 ( .IN1(n30), .IN2(\data_i[1][7] ), .IN3(n14), .IN4(
        \data_i[0][7] ), .Q(n637) );
  AO22X1 U667 ( .IN1(n31), .IN2(\data_i[6][7] ), .IN3(n15), .IN4(
        \data_i[7][7] ), .Q(n636) );
  AO22X1 U668 ( .IN1(n32), .IN2(\data_i[5][7] ), .IN3(n16), .IN4(
        \data_i[4][7] ), .Q(n635) );
  NOR4X0 U669 ( .IN1(n638), .IN2(n637), .IN3(n636), .IN4(n635), .QN(n649) );
  AO22X1 U670 ( .IN1(n17), .IN2(\data_i[26][7] ), .IN3(n1), .IN4(
        \data_i[27][7] ), .Q(n642) );
  AO22X1 U671 ( .IN1(n18), .IN2(\data_i[25][7] ), .IN3(n2), .IN4(
        \data_i[24][7] ), .Q(n641) );
  AO22X1 U672 ( .IN1(n19), .IN2(\data_i[30][7] ), .IN3(n3), .IN4(
        \data_i[31][7] ), .Q(n640) );
  AO22X1 U673 ( .IN1(n20), .IN2(\data_i[29][7] ), .IN3(n4), .IN4(
        \data_i[28][7] ), .Q(n639) );
  NOR4X0 U674 ( .IN1(n642), .IN2(n641), .IN3(n640), .IN4(n639), .QN(n648) );
  AO22X1 U675 ( .IN1(n21), .IN2(\data_i[18][7] ), .IN3(n5), .IN4(
        \data_i[19][7] ), .Q(n646) );
  AO22X1 U676 ( .IN1(n22), .IN2(\data_i[17][7] ), .IN3(n6), .IN4(
        \data_i[16][7] ), .Q(n645) );
  AO22X1 U677 ( .IN1(n23), .IN2(\data_i[22][7] ), .IN3(n7), .IN4(
        \data_i[23][7] ), .Q(n644) );
  AO22X1 U678 ( .IN1(n24), .IN2(\data_i[21][7] ), .IN3(n8), .IN4(
        \data_i[20][7] ), .Q(n643) );
  NOR4X0 U679 ( .IN1(n646), .IN2(n645), .IN3(n644), .IN4(n643), .QN(n647) );
  NAND4X0 U680 ( .IN1(n650), .IN2(n649), .IN3(n648), .IN4(n647), .QN(data_o[7]) );
  AO22X1 U681 ( .IN1(n25), .IN2(\data_i[10][8] ), .IN3(n9), .IN4(
        \data_i[11][8] ), .Q(n654) );
  AO22X1 U682 ( .IN1(n26), .IN2(\data_i[9][8] ), .IN3(n10), .IN4(
        \data_i[8][8] ), .Q(n653) );
  AO22X1 U683 ( .IN1(n27), .IN2(\data_i[14][8] ), .IN3(n11), .IN4(
        \data_i[15][8] ), .Q(n652) );
  AO22X1 U684 ( .IN1(n28), .IN2(\data_i[13][8] ), .IN3(n12), .IN4(
        \data_i[12][8] ), .Q(n651) );
  NOR4X0 U685 ( .IN1(n654), .IN2(n653), .IN3(n652), .IN4(n651), .QN(n670) );
  AO22X1 U686 ( .IN1(n29), .IN2(\data_i[2][8] ), .IN3(n13), .IN4(
        \data_i[3][8] ), .Q(n658) );
  AO22X1 U687 ( .IN1(n30), .IN2(\data_i[1][8] ), .IN3(n14), .IN4(
        \data_i[0][8] ), .Q(n657) );
  AO22X1 U688 ( .IN1(n31), .IN2(\data_i[6][8] ), .IN3(n15), .IN4(
        \data_i[7][8] ), .Q(n656) );
  AO22X1 U689 ( .IN1(n32), .IN2(\data_i[5][8] ), .IN3(n16), .IN4(
        \data_i[4][8] ), .Q(n655) );
  NOR4X0 U690 ( .IN1(n658), .IN2(n657), .IN3(n656), .IN4(n655), .QN(n669) );
  AO22X1 U691 ( .IN1(n17), .IN2(\data_i[26][8] ), .IN3(n1), .IN4(
        \data_i[27][8] ), .Q(n662) );
  AO22X1 U692 ( .IN1(n18), .IN2(\data_i[25][8] ), .IN3(n2), .IN4(
        \data_i[24][8] ), .Q(n661) );
  AO22X1 U693 ( .IN1(n19), .IN2(\data_i[30][8] ), .IN3(n3), .IN4(
        \data_i[31][8] ), .Q(n660) );
  AO22X1 U694 ( .IN1(n20), .IN2(\data_i[29][8] ), .IN3(n4), .IN4(
        \data_i[28][8] ), .Q(n659) );
  NOR4X0 U695 ( .IN1(n662), .IN2(n661), .IN3(n660), .IN4(n659), .QN(n668) );
  AO22X1 U696 ( .IN1(n21), .IN2(\data_i[18][8] ), .IN3(n5), .IN4(
        \data_i[19][8] ), .Q(n666) );
  AO22X1 U697 ( .IN1(n22), .IN2(\data_i[17][8] ), .IN3(n6), .IN4(
        \data_i[16][8] ), .Q(n665) );
  AO22X1 U698 ( .IN1(n23), .IN2(\data_i[22][8] ), .IN3(n7), .IN4(
        \data_i[23][8] ), .Q(n664) );
  AO22X1 U699 ( .IN1(n24), .IN2(\data_i[21][8] ), .IN3(n8), .IN4(
        \data_i[20][8] ), .Q(n663) );
  NOR4X0 U700 ( .IN1(n666), .IN2(n665), .IN3(n664), .IN4(n663), .QN(n667) );
  NAND4X0 U701 ( .IN1(n670), .IN2(n669), .IN3(n668), .IN4(n667), .QN(data_o[8]) );
  AO22X1 U702 ( .IN1(n25), .IN2(\data_i[10][9] ), .IN3(n9), .IN4(
        \data_i[11][9] ), .Q(n674) );
  AO22X1 U703 ( .IN1(n26), .IN2(\data_i[9][9] ), .IN3(n10), .IN4(
        \data_i[8][9] ), .Q(n673) );
  AO22X1 U704 ( .IN1(n27), .IN2(\data_i[14][9] ), .IN3(n11), .IN4(
        \data_i[15][9] ), .Q(n672) );
  AO22X1 U705 ( .IN1(n28), .IN2(\data_i[13][9] ), .IN3(n12), .IN4(
        \data_i[12][9] ), .Q(n671) );
  NOR4X0 U706 ( .IN1(n674), .IN2(n673), .IN3(n672), .IN4(n671), .QN(n690) );
  AO22X1 U707 ( .IN1(n29), .IN2(\data_i[2][9] ), .IN3(n13), .IN4(
        \data_i[3][9] ), .Q(n678) );
  AO22X1 U708 ( .IN1(n30), .IN2(\data_i[1][9] ), .IN3(n14), .IN4(
        \data_i[0][9] ), .Q(n677) );
  AO22X1 U709 ( .IN1(n31), .IN2(\data_i[6][9] ), .IN3(n15), .IN4(
        \data_i[7][9] ), .Q(n676) );
  AO22X1 U710 ( .IN1(n32), .IN2(\data_i[5][9] ), .IN3(n16), .IN4(
        \data_i[4][9] ), .Q(n675) );
  NOR4X0 U711 ( .IN1(n678), .IN2(n677), .IN3(n676), .IN4(n675), .QN(n689) );
  AO22X1 U712 ( .IN1(n17), .IN2(\data_i[26][9] ), .IN3(n1), .IN4(
        \data_i[27][9] ), .Q(n682) );
  AO22X1 U713 ( .IN1(n18), .IN2(\data_i[25][9] ), .IN3(n2), .IN4(
        \data_i[24][9] ), .Q(n681) );
  AO22X1 U714 ( .IN1(n19), .IN2(\data_i[30][9] ), .IN3(n3), .IN4(
        \data_i[31][9] ), .Q(n680) );
  AO22X1 U715 ( .IN1(n20), .IN2(\data_i[29][9] ), .IN3(n4), .IN4(
        \data_i[28][9] ), .Q(n679) );
  NOR4X0 U716 ( .IN1(n682), .IN2(n681), .IN3(n680), .IN4(n679), .QN(n688) );
  AO22X1 U717 ( .IN1(n21), .IN2(\data_i[18][9] ), .IN3(n5), .IN4(
        \data_i[19][9] ), .Q(n686) );
  AO22X1 U718 ( .IN1(n22), .IN2(\data_i[17][9] ), .IN3(n6), .IN4(
        \data_i[16][9] ), .Q(n685) );
  AO22X1 U719 ( .IN1(n23), .IN2(\data_i[22][9] ), .IN3(n7), .IN4(
        \data_i[23][9] ), .Q(n684) );
  AO22X1 U720 ( .IN1(n24), .IN2(\data_i[21][9] ), .IN3(n8), .IN4(
        \data_i[20][9] ), .Q(n683) );
  NOR4X0 U721 ( .IN1(n686), .IN2(n685), .IN3(n684), .IN4(n683), .QN(n687) );
  NAND4X0 U722 ( .IN1(n690), .IN2(n689), .IN3(n688), .IN4(n687), .QN(data_o[9]) );
endmodule


module cam ( reset, clk, read, read_index, write, write_index, write_data, 
        search, search_data, read_valid, read_value, search_valid, 
        search_index );
  input [4:0] read_index;
  input [4:0] write_index;
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  output [4:0] search_index;
  input reset, clk, read, write, search;
  output read_valid, search_valid;
  wire   \read_value_mux[31][31] , \read_value_mux[31][30] ,
         \read_value_mux[31][29] , \read_value_mux[31][28] ,
         \read_value_mux[31][27] , \read_value_mux[31][26] ,
         \read_value_mux[31][25] , \read_value_mux[31][24] ,
         \read_value_mux[31][23] , \read_value_mux[31][22] ,
         \read_value_mux[31][21] , \read_value_mux[31][20] ,
         \read_value_mux[31][19] , \read_value_mux[31][18] ,
         \read_value_mux[31][17] , \read_value_mux[31][16] ,
         \read_value_mux[31][15] , \read_value_mux[31][14] ,
         \read_value_mux[31][13] , \read_value_mux[31][12] ,
         \read_value_mux[31][11] , \read_value_mux[31][10] ,
         \read_value_mux[31][9] , \read_value_mux[31][8] ,
         \read_value_mux[31][7] , \read_value_mux[31][6] ,
         \read_value_mux[31][5] , \read_value_mux[31][4] ,
         \read_value_mux[31][3] , \read_value_mux[31][2] ,
         \read_value_mux[31][1] , \read_value_mux[31][0] ,
         \read_value_mux[30][31] , \read_value_mux[30][30] ,
         \read_value_mux[30][29] , \read_value_mux[30][28] ,
         \read_value_mux[30][27] , \read_value_mux[30][26] ,
         \read_value_mux[30][25] , \read_value_mux[30][24] ,
         \read_value_mux[30][23] , \read_value_mux[30][22] ,
         \read_value_mux[30][21] , \read_value_mux[30][20] ,
         \read_value_mux[30][19] , \read_value_mux[30][18] ,
         \read_value_mux[30][17] , \read_value_mux[30][16] ,
         \read_value_mux[30][15] , \read_value_mux[30][14] ,
         \read_value_mux[30][13] , \read_value_mux[30][12] ,
         \read_value_mux[30][11] , \read_value_mux[30][10] ,
         \read_value_mux[30][9] , \read_value_mux[30][8] ,
         \read_value_mux[30][7] , \read_value_mux[30][6] ,
         \read_value_mux[30][5] , \read_value_mux[30][4] ,
         \read_value_mux[30][3] , \read_value_mux[30][2] ,
         \read_value_mux[30][1] , \read_value_mux[30][0] ,
         \read_value_mux[29][31] , \read_value_mux[29][30] ,
         \read_value_mux[29][29] , \read_value_mux[29][28] ,
         \read_value_mux[29][27] , \read_value_mux[29][26] ,
         \read_value_mux[29][25] , \read_value_mux[29][24] ,
         \read_value_mux[29][23] , \read_value_mux[29][22] ,
         \read_value_mux[29][21] , \read_value_mux[29][20] ,
         \read_value_mux[29][19] , \read_value_mux[29][18] ,
         \read_value_mux[29][17] , \read_value_mux[29][16] ,
         \read_value_mux[29][15] , \read_value_mux[29][14] ,
         \read_value_mux[29][13] , \read_value_mux[29][12] ,
         \read_value_mux[29][11] , \read_value_mux[29][10] ,
         \read_value_mux[29][9] , \read_value_mux[29][8] ,
         \read_value_mux[29][7] , \read_value_mux[29][6] ,
         \read_value_mux[29][5] , \read_value_mux[29][4] ,
         \read_value_mux[29][3] , \read_value_mux[29][2] ,
         \read_value_mux[29][1] , \read_value_mux[29][0] ,
         \read_value_mux[28][31] , \read_value_mux[28][30] ,
         \read_value_mux[28][29] , \read_value_mux[28][28] ,
         \read_value_mux[28][27] , \read_value_mux[28][26] ,
         \read_value_mux[28][25] , \read_value_mux[28][24] ,
         \read_value_mux[28][23] , \read_value_mux[28][22] ,
         \read_value_mux[28][21] , \read_value_mux[28][20] ,
         \read_value_mux[28][19] , \read_value_mux[28][18] ,
         \read_value_mux[28][17] , \read_value_mux[28][16] ,
         \read_value_mux[28][15] , \read_value_mux[28][14] ,
         \read_value_mux[28][13] , \read_value_mux[28][12] ,
         \read_value_mux[28][11] , \read_value_mux[28][10] ,
         \read_value_mux[28][9] , \read_value_mux[28][8] ,
         \read_value_mux[28][7] , \read_value_mux[28][6] ,
         \read_value_mux[28][5] , \read_value_mux[28][4] ,
         \read_value_mux[28][3] , \read_value_mux[28][2] ,
         \read_value_mux[28][1] , \read_value_mux[28][0] ,
         \read_value_mux[27][31] , \read_value_mux[27][30] ,
         \read_value_mux[27][29] , \read_value_mux[27][28] ,
         \read_value_mux[27][27] , \read_value_mux[27][26] ,
         \read_value_mux[27][25] , \read_value_mux[27][24] ,
         \read_value_mux[27][23] , \read_value_mux[27][22] ,
         \read_value_mux[27][21] , \read_value_mux[27][20] ,
         \read_value_mux[27][19] , \read_value_mux[27][18] ,
         \read_value_mux[27][17] , \read_value_mux[27][16] ,
         \read_value_mux[27][15] , \read_value_mux[27][14] ,
         \read_value_mux[27][13] , \read_value_mux[27][12] ,
         \read_value_mux[27][11] , \read_value_mux[27][10] ,
         \read_value_mux[27][9] , \read_value_mux[27][8] ,
         \read_value_mux[27][7] , \read_value_mux[27][6] ,
         \read_value_mux[27][5] , \read_value_mux[27][4] ,
         \read_value_mux[27][3] , \read_value_mux[27][2] ,
         \read_value_mux[27][1] , \read_value_mux[27][0] ,
         \read_value_mux[26][31] , \read_value_mux[26][30] ,
         \read_value_mux[26][29] , \read_value_mux[26][28] ,
         \read_value_mux[26][27] , \read_value_mux[26][26] ,
         \read_value_mux[26][25] , \read_value_mux[26][24] ,
         \read_value_mux[26][23] , \read_value_mux[26][22] ,
         \read_value_mux[26][21] , \read_value_mux[26][20] ,
         \read_value_mux[26][19] , \read_value_mux[26][18] ,
         \read_value_mux[26][17] , \read_value_mux[26][16] ,
         \read_value_mux[26][15] , \read_value_mux[26][14] ,
         \read_value_mux[26][13] , \read_value_mux[26][12] ,
         \read_value_mux[26][11] , \read_value_mux[26][10] ,
         \read_value_mux[26][9] , \read_value_mux[26][8] ,
         \read_value_mux[26][7] , \read_value_mux[26][6] ,
         \read_value_mux[26][5] , \read_value_mux[26][4] ,
         \read_value_mux[26][3] , \read_value_mux[26][2] ,
         \read_value_mux[26][1] , \read_value_mux[26][0] ,
         \read_value_mux[25][31] , \read_value_mux[25][30] ,
         \read_value_mux[25][29] , \read_value_mux[25][28] ,
         \read_value_mux[25][27] , \read_value_mux[25][26] ,
         \read_value_mux[25][25] , \read_value_mux[25][24] ,
         \read_value_mux[25][23] , \read_value_mux[25][22] ,
         \read_value_mux[25][21] , \read_value_mux[25][20] ,
         \read_value_mux[25][19] , \read_value_mux[25][18] ,
         \read_value_mux[25][17] , \read_value_mux[25][16] ,
         \read_value_mux[25][15] , \read_value_mux[25][14] ,
         \read_value_mux[25][13] , \read_value_mux[25][12] ,
         \read_value_mux[25][11] , \read_value_mux[25][10] ,
         \read_value_mux[25][9] , \read_value_mux[25][8] ,
         \read_value_mux[25][7] , \read_value_mux[25][6] ,
         \read_value_mux[25][5] , \read_value_mux[25][4] ,
         \read_value_mux[25][3] , \read_value_mux[25][2] ,
         \read_value_mux[25][1] , \read_value_mux[25][0] ,
         \read_value_mux[24][31] , \read_value_mux[24][30] ,
         \read_value_mux[24][29] , \read_value_mux[24][28] ,
         \read_value_mux[24][27] , \read_value_mux[24][26] ,
         \read_value_mux[24][25] , \read_value_mux[24][24] ,
         \read_value_mux[24][23] , \read_value_mux[24][22] ,
         \read_value_mux[24][21] , \read_value_mux[24][20] ,
         \read_value_mux[24][19] , \read_value_mux[24][18] ,
         \read_value_mux[24][17] , \read_value_mux[24][16] ,
         \read_value_mux[24][15] , \read_value_mux[24][14] ,
         \read_value_mux[24][13] , \read_value_mux[24][12] ,
         \read_value_mux[24][11] , \read_value_mux[24][10] ,
         \read_value_mux[24][9] , \read_value_mux[24][8] ,
         \read_value_mux[24][7] , \read_value_mux[24][6] ,
         \read_value_mux[24][5] , \read_value_mux[24][4] ,
         \read_value_mux[24][3] , \read_value_mux[24][2] ,
         \read_value_mux[24][1] , \read_value_mux[24][0] ,
         \read_value_mux[23][31] , \read_value_mux[23][30] ,
         \read_value_mux[23][29] , \read_value_mux[23][28] ,
         \read_value_mux[23][27] , \read_value_mux[23][26] ,
         \read_value_mux[23][25] , \read_value_mux[23][24] ,
         \read_value_mux[23][23] , \read_value_mux[23][22] ,
         \read_value_mux[23][21] , \read_value_mux[23][20] ,
         \read_value_mux[23][19] , \read_value_mux[23][18] ,
         \read_value_mux[23][17] , \read_value_mux[23][16] ,
         \read_value_mux[23][15] , \read_value_mux[23][14] ,
         \read_value_mux[23][13] , \read_value_mux[23][12] ,
         \read_value_mux[23][11] , \read_value_mux[23][10] ,
         \read_value_mux[23][9] , \read_value_mux[23][8] ,
         \read_value_mux[23][7] , \read_value_mux[23][6] ,
         \read_value_mux[23][5] , \read_value_mux[23][4] ,
         \read_value_mux[23][3] , \read_value_mux[23][2] ,
         \read_value_mux[23][1] , \read_value_mux[23][0] ,
         \read_value_mux[22][31] , \read_value_mux[22][30] ,
         \read_value_mux[22][29] , \read_value_mux[22][28] ,
         \read_value_mux[22][27] , \read_value_mux[22][26] ,
         \read_value_mux[22][25] , \read_value_mux[22][24] ,
         \read_value_mux[22][23] , \read_value_mux[22][22] ,
         \read_value_mux[22][21] , \read_value_mux[22][20] ,
         \read_value_mux[22][19] , \read_value_mux[22][18] ,
         \read_value_mux[22][17] , \read_value_mux[22][16] ,
         \read_value_mux[22][15] , \read_value_mux[22][14] ,
         \read_value_mux[22][13] , \read_value_mux[22][12] ,
         \read_value_mux[22][11] , \read_value_mux[22][10] ,
         \read_value_mux[22][9] , \read_value_mux[22][8] ,
         \read_value_mux[22][7] , \read_value_mux[22][6] ,
         \read_value_mux[22][5] , \read_value_mux[22][4] ,
         \read_value_mux[22][3] , \read_value_mux[22][2] ,
         \read_value_mux[22][1] , \read_value_mux[22][0] ,
         \read_value_mux[21][31] , \read_value_mux[21][30] ,
         \read_value_mux[21][29] , \read_value_mux[21][28] ,
         \read_value_mux[21][27] , \read_value_mux[21][26] ,
         \read_value_mux[21][25] , \read_value_mux[21][24] ,
         \read_value_mux[21][23] , \read_value_mux[21][22] ,
         \read_value_mux[21][21] , \read_value_mux[21][20] ,
         \read_value_mux[21][19] , \read_value_mux[21][18] ,
         \read_value_mux[21][17] , \read_value_mux[21][16] ,
         \read_value_mux[21][15] , \read_value_mux[21][14] ,
         \read_value_mux[21][13] , \read_value_mux[21][12] ,
         \read_value_mux[21][11] , \read_value_mux[21][10] ,
         \read_value_mux[21][9] , \read_value_mux[21][8] ,
         \read_value_mux[21][7] , \read_value_mux[21][6] ,
         \read_value_mux[21][5] , \read_value_mux[21][4] ,
         \read_value_mux[21][3] , \read_value_mux[21][2] ,
         \read_value_mux[21][1] , \read_value_mux[21][0] ,
         \read_value_mux[20][31] , \read_value_mux[20][30] ,
         \read_value_mux[20][29] , \read_value_mux[20][28] ,
         \read_value_mux[20][27] , \read_value_mux[20][26] ,
         \read_value_mux[20][25] , \read_value_mux[20][24] ,
         \read_value_mux[20][23] , \read_value_mux[20][22] ,
         \read_value_mux[20][21] , \read_value_mux[20][20] ,
         \read_value_mux[20][19] , \read_value_mux[20][18] ,
         \read_value_mux[20][17] , \read_value_mux[20][16] ,
         \read_value_mux[20][15] , \read_value_mux[20][14] ,
         \read_value_mux[20][13] , \read_value_mux[20][12] ,
         \read_value_mux[20][11] , \read_value_mux[20][10] ,
         \read_value_mux[20][9] , \read_value_mux[20][8] ,
         \read_value_mux[20][7] , \read_value_mux[20][6] ,
         \read_value_mux[20][5] , \read_value_mux[20][4] ,
         \read_value_mux[20][3] , \read_value_mux[20][2] ,
         \read_value_mux[20][1] , \read_value_mux[20][0] ,
         \read_value_mux[19][31] , \read_value_mux[19][30] ,
         \read_value_mux[19][29] , \read_value_mux[19][28] ,
         \read_value_mux[19][27] , \read_value_mux[19][26] ,
         \read_value_mux[19][25] , \read_value_mux[19][24] ,
         \read_value_mux[19][23] , \read_value_mux[19][22] ,
         \read_value_mux[19][21] , \read_value_mux[19][20] ,
         \read_value_mux[19][19] , \read_value_mux[19][18] ,
         \read_value_mux[19][17] , \read_value_mux[19][16] ,
         \read_value_mux[19][15] , \read_value_mux[19][14] ,
         \read_value_mux[19][13] , \read_value_mux[19][12] ,
         \read_value_mux[19][11] , \read_value_mux[19][10] ,
         \read_value_mux[19][9] , \read_value_mux[19][8] ,
         \read_value_mux[19][7] , \read_value_mux[19][6] ,
         \read_value_mux[19][5] , \read_value_mux[19][4] ,
         \read_value_mux[19][3] , \read_value_mux[19][2] ,
         \read_value_mux[19][1] , \read_value_mux[19][0] ,
         \read_value_mux[18][31] , \read_value_mux[18][30] ,
         \read_value_mux[18][29] , \read_value_mux[18][28] ,
         \read_value_mux[18][27] , \read_value_mux[18][26] ,
         \read_value_mux[18][25] , \read_value_mux[18][24] ,
         \read_value_mux[18][23] , \read_value_mux[18][22] ,
         \read_value_mux[18][21] , \read_value_mux[18][20] ,
         \read_value_mux[18][19] , \read_value_mux[18][18] ,
         \read_value_mux[18][17] , \read_value_mux[18][16] ,
         \read_value_mux[18][15] , \read_value_mux[18][14] ,
         \read_value_mux[18][13] , \read_value_mux[18][12] ,
         \read_value_mux[18][11] , \read_value_mux[18][10] ,
         \read_value_mux[18][9] , \read_value_mux[18][8] ,
         \read_value_mux[18][7] , \read_value_mux[18][6] ,
         \read_value_mux[18][5] , \read_value_mux[18][4] ,
         \read_value_mux[18][3] , \read_value_mux[18][2] ,
         \read_value_mux[18][1] , \read_value_mux[18][0] ,
         \read_value_mux[17][31] , \read_value_mux[17][30] ,
         \read_value_mux[17][29] , \read_value_mux[17][28] ,
         \read_value_mux[17][27] , \read_value_mux[17][26] ,
         \read_value_mux[17][25] , \read_value_mux[17][24] ,
         \read_value_mux[17][23] , \read_value_mux[17][22] ,
         \read_value_mux[17][21] , \read_value_mux[17][20] ,
         \read_value_mux[17][19] , \read_value_mux[17][18] ,
         \read_value_mux[17][17] , \read_value_mux[17][16] ,
         \read_value_mux[17][15] , \read_value_mux[17][14] ,
         \read_value_mux[17][13] , \read_value_mux[17][12] ,
         \read_value_mux[17][11] , \read_value_mux[17][10] ,
         \read_value_mux[17][9] , \read_value_mux[17][8] ,
         \read_value_mux[17][7] , \read_value_mux[17][6] ,
         \read_value_mux[17][5] , \read_value_mux[17][4] ,
         \read_value_mux[17][3] , \read_value_mux[17][2] ,
         \read_value_mux[17][1] , \read_value_mux[17][0] ,
         \read_value_mux[16][31] , \read_value_mux[16][30] ,
         \read_value_mux[16][29] , \read_value_mux[16][28] ,
         \read_value_mux[16][27] , \read_value_mux[16][26] ,
         \read_value_mux[16][25] , \read_value_mux[16][24] ,
         \read_value_mux[16][23] , \read_value_mux[16][22] ,
         \read_value_mux[16][21] , \read_value_mux[16][20] ,
         \read_value_mux[16][19] , \read_value_mux[16][18] ,
         \read_value_mux[16][17] , \read_value_mux[16][16] ,
         \read_value_mux[16][15] , \read_value_mux[16][14] ,
         \read_value_mux[16][13] , \read_value_mux[16][12] ,
         \read_value_mux[16][11] , \read_value_mux[16][10] ,
         \read_value_mux[16][9] , \read_value_mux[16][8] ,
         \read_value_mux[16][7] , \read_value_mux[16][6] ,
         \read_value_mux[16][5] , \read_value_mux[16][4] ,
         \read_value_mux[16][3] , \read_value_mux[16][2] ,
         \read_value_mux[16][1] , \read_value_mux[16][0] ,
         \read_value_mux[15][31] , \read_value_mux[15][30] ,
         \read_value_mux[15][29] , \read_value_mux[15][28] ,
         \read_value_mux[15][27] , \read_value_mux[15][26] ,
         \read_value_mux[15][25] , \read_value_mux[15][24] ,
         \read_value_mux[15][23] , \read_value_mux[15][22] ,
         \read_value_mux[15][21] , \read_value_mux[15][20] ,
         \read_value_mux[15][19] , \read_value_mux[15][18] ,
         \read_value_mux[15][17] , \read_value_mux[15][16] ,
         \read_value_mux[15][15] , \read_value_mux[15][14] ,
         \read_value_mux[15][13] , \read_value_mux[15][12] ,
         \read_value_mux[15][11] , \read_value_mux[15][10] ,
         \read_value_mux[15][9] , \read_value_mux[15][8] ,
         \read_value_mux[15][7] , \read_value_mux[15][6] ,
         \read_value_mux[15][5] , \read_value_mux[15][4] ,
         \read_value_mux[15][3] , \read_value_mux[15][2] ,
         \read_value_mux[15][1] , \read_value_mux[15][0] ,
         \read_value_mux[14][31] , \read_value_mux[14][30] ,
         \read_value_mux[14][29] , \read_value_mux[14][28] ,
         \read_value_mux[14][27] , \read_value_mux[14][26] ,
         \read_value_mux[14][25] , \read_value_mux[14][24] ,
         \read_value_mux[14][23] , \read_value_mux[14][22] ,
         \read_value_mux[14][21] , \read_value_mux[14][20] ,
         \read_value_mux[14][19] , \read_value_mux[14][18] ,
         \read_value_mux[14][17] , \read_value_mux[14][16] ,
         \read_value_mux[14][15] , \read_value_mux[14][14] ,
         \read_value_mux[14][13] , \read_value_mux[14][12] ,
         \read_value_mux[14][11] , \read_value_mux[14][10] ,
         \read_value_mux[14][9] , \read_value_mux[14][8] ,
         \read_value_mux[14][7] , \read_value_mux[14][6] ,
         \read_value_mux[14][5] , \read_value_mux[14][4] ,
         \read_value_mux[14][3] , \read_value_mux[14][2] ,
         \read_value_mux[14][1] , \read_value_mux[14][0] ,
         \read_value_mux[13][31] , \read_value_mux[13][30] ,
         \read_value_mux[13][29] , \read_value_mux[13][28] ,
         \read_value_mux[13][27] , \read_value_mux[13][26] ,
         \read_value_mux[13][25] , \read_value_mux[13][24] ,
         \read_value_mux[13][23] , \read_value_mux[13][22] ,
         \read_value_mux[13][21] , \read_value_mux[13][20] ,
         \read_value_mux[13][19] , \read_value_mux[13][18] ,
         \read_value_mux[13][17] , \read_value_mux[13][16] ,
         \read_value_mux[13][15] , \read_value_mux[13][14] ,
         \read_value_mux[13][13] , \read_value_mux[13][12] ,
         \read_value_mux[13][11] , \read_value_mux[13][10] ,
         \read_value_mux[13][9] , \read_value_mux[13][8] ,
         \read_value_mux[13][7] , \read_value_mux[13][6] ,
         \read_value_mux[13][5] , \read_value_mux[13][4] ,
         \read_value_mux[13][3] , \read_value_mux[13][2] ,
         \read_value_mux[13][1] , \read_value_mux[13][0] ,
         \read_value_mux[12][31] , \read_value_mux[12][30] ,
         \read_value_mux[12][29] , \read_value_mux[12][28] ,
         \read_value_mux[12][27] , \read_value_mux[12][26] ,
         \read_value_mux[12][25] , \read_value_mux[12][24] ,
         \read_value_mux[12][23] , \read_value_mux[12][22] ,
         \read_value_mux[12][21] , \read_value_mux[12][20] ,
         \read_value_mux[12][19] , \read_value_mux[12][18] ,
         \read_value_mux[12][17] , \read_value_mux[12][16] ,
         \read_value_mux[12][15] , \read_value_mux[12][14] ,
         \read_value_mux[12][13] , \read_value_mux[12][12] ,
         \read_value_mux[12][11] , \read_value_mux[12][10] ,
         \read_value_mux[12][9] , \read_value_mux[12][8] ,
         \read_value_mux[12][7] , \read_value_mux[12][6] ,
         \read_value_mux[12][5] , \read_value_mux[12][4] ,
         \read_value_mux[12][3] , \read_value_mux[12][2] ,
         \read_value_mux[12][1] , \read_value_mux[12][0] ,
         \read_value_mux[11][31] , \read_value_mux[11][30] ,
         \read_value_mux[11][29] , \read_value_mux[11][28] ,
         \read_value_mux[11][27] , \read_value_mux[11][26] ,
         \read_value_mux[11][25] , \read_value_mux[11][24] ,
         \read_value_mux[11][23] , \read_value_mux[11][22] ,
         \read_value_mux[11][21] , \read_value_mux[11][20] ,
         \read_value_mux[11][19] , \read_value_mux[11][18] ,
         \read_value_mux[11][17] , \read_value_mux[11][16] ,
         \read_value_mux[11][15] , \read_value_mux[11][14] ,
         \read_value_mux[11][13] , \read_value_mux[11][12] ,
         \read_value_mux[11][11] , \read_value_mux[11][10] ,
         \read_value_mux[11][9] , \read_value_mux[11][8] ,
         \read_value_mux[11][7] , \read_value_mux[11][6] ,
         \read_value_mux[11][5] , \read_value_mux[11][4] ,
         \read_value_mux[11][3] , \read_value_mux[11][2] ,
         \read_value_mux[11][1] , \read_value_mux[11][0] ,
         \read_value_mux[10][31] , \read_value_mux[10][30] ,
         \read_value_mux[10][29] , \read_value_mux[10][28] ,
         \read_value_mux[10][27] , \read_value_mux[10][26] ,
         \read_value_mux[10][25] , \read_value_mux[10][24] ,
         \read_value_mux[10][23] , \read_value_mux[10][22] ,
         \read_value_mux[10][21] , \read_value_mux[10][20] ,
         \read_value_mux[10][19] , \read_value_mux[10][18] ,
         \read_value_mux[10][17] , \read_value_mux[10][16] ,
         \read_value_mux[10][15] , \read_value_mux[10][14] ,
         \read_value_mux[10][13] , \read_value_mux[10][12] ,
         \read_value_mux[10][11] , \read_value_mux[10][10] ,
         \read_value_mux[10][9] , \read_value_mux[10][8] ,
         \read_value_mux[10][7] , \read_value_mux[10][6] ,
         \read_value_mux[10][5] , \read_value_mux[10][4] ,
         \read_value_mux[10][3] , \read_value_mux[10][2] ,
         \read_value_mux[10][1] , \read_value_mux[10][0] ,
         \read_value_mux[9][31] , \read_value_mux[9][30] ,
         \read_value_mux[9][29] , \read_value_mux[9][28] ,
         \read_value_mux[9][27] , \read_value_mux[9][26] ,
         \read_value_mux[9][25] , \read_value_mux[9][24] ,
         \read_value_mux[9][23] , \read_value_mux[9][22] ,
         \read_value_mux[9][21] , \read_value_mux[9][20] ,
         \read_value_mux[9][19] , \read_value_mux[9][18] ,
         \read_value_mux[9][17] , \read_value_mux[9][16] ,
         \read_value_mux[9][15] , \read_value_mux[9][14] ,
         \read_value_mux[9][13] , \read_value_mux[9][12] ,
         \read_value_mux[9][11] , \read_value_mux[9][10] ,
         \read_value_mux[9][9] , \read_value_mux[9][8] ,
         \read_value_mux[9][7] , \read_value_mux[9][6] ,
         \read_value_mux[9][5] , \read_value_mux[9][4] ,
         \read_value_mux[9][3] , \read_value_mux[9][2] ,
         \read_value_mux[9][1] , \read_value_mux[9][0] ,
         \read_value_mux[8][31] , \read_value_mux[8][30] ,
         \read_value_mux[8][29] , \read_value_mux[8][28] ,
         \read_value_mux[8][27] , \read_value_mux[8][26] ,
         \read_value_mux[8][25] , \read_value_mux[8][24] ,
         \read_value_mux[8][23] , \read_value_mux[8][22] ,
         \read_value_mux[8][21] , \read_value_mux[8][20] ,
         \read_value_mux[8][19] , \read_value_mux[8][18] ,
         \read_value_mux[8][17] , \read_value_mux[8][16] ,
         \read_value_mux[8][15] , \read_value_mux[8][14] ,
         \read_value_mux[8][13] , \read_value_mux[8][12] ,
         \read_value_mux[8][11] , \read_value_mux[8][10] ,
         \read_value_mux[8][9] , \read_value_mux[8][8] ,
         \read_value_mux[8][7] , \read_value_mux[8][6] ,
         \read_value_mux[8][5] , \read_value_mux[8][4] ,
         \read_value_mux[8][3] , \read_value_mux[8][2] ,
         \read_value_mux[8][1] , \read_value_mux[8][0] ,
         \read_value_mux[7][31] , \read_value_mux[7][30] ,
         \read_value_mux[7][29] , \read_value_mux[7][28] ,
         \read_value_mux[7][27] , \read_value_mux[7][26] ,
         \read_value_mux[7][25] , \read_value_mux[7][24] ,
         \read_value_mux[7][23] , \read_value_mux[7][22] ,
         \read_value_mux[7][21] , \read_value_mux[7][20] ,
         \read_value_mux[7][19] , \read_value_mux[7][18] ,
         \read_value_mux[7][17] , \read_value_mux[7][16] ,
         \read_value_mux[7][15] , \read_value_mux[7][14] ,
         \read_value_mux[7][13] , \read_value_mux[7][12] ,
         \read_value_mux[7][11] , \read_value_mux[7][10] ,
         \read_value_mux[7][9] , \read_value_mux[7][8] ,
         \read_value_mux[7][7] , \read_value_mux[7][6] ,
         \read_value_mux[7][5] , \read_value_mux[7][4] ,
         \read_value_mux[7][3] , \read_value_mux[7][2] ,
         \read_value_mux[7][1] , \read_value_mux[7][0] ,
         \read_value_mux[6][31] , \read_value_mux[6][30] ,
         \read_value_mux[6][29] , \read_value_mux[6][28] ,
         \read_value_mux[6][27] , \read_value_mux[6][26] ,
         \read_value_mux[6][25] , \read_value_mux[6][24] ,
         \read_value_mux[6][23] , \read_value_mux[6][22] ,
         \read_value_mux[6][21] , \read_value_mux[6][20] ,
         \read_value_mux[6][19] , \read_value_mux[6][18] ,
         \read_value_mux[6][17] , \read_value_mux[6][16] ,
         \read_value_mux[6][15] , \read_value_mux[6][14] ,
         \read_value_mux[6][13] , \read_value_mux[6][12] ,
         \read_value_mux[6][11] , \read_value_mux[6][10] ,
         \read_value_mux[6][9] , \read_value_mux[6][8] ,
         \read_value_mux[6][7] , \read_value_mux[6][6] ,
         \read_value_mux[6][5] , \read_value_mux[6][4] ,
         \read_value_mux[6][3] , \read_value_mux[6][2] ,
         \read_value_mux[6][1] , \read_value_mux[6][0] ,
         \read_value_mux[5][31] , \read_value_mux[5][30] ,
         \read_value_mux[5][29] , \read_value_mux[5][28] ,
         \read_value_mux[5][27] , \read_value_mux[5][26] ,
         \read_value_mux[5][25] , \read_value_mux[5][24] ,
         \read_value_mux[5][23] , \read_value_mux[5][22] ,
         \read_value_mux[5][21] , \read_value_mux[5][20] ,
         \read_value_mux[5][19] , \read_value_mux[5][18] ,
         \read_value_mux[5][17] , \read_value_mux[5][16] ,
         \read_value_mux[5][15] , \read_value_mux[5][14] ,
         \read_value_mux[5][13] , \read_value_mux[5][12] ,
         \read_value_mux[5][11] , \read_value_mux[5][10] ,
         \read_value_mux[5][9] , \read_value_mux[5][8] ,
         \read_value_mux[5][7] , \read_value_mux[5][6] ,
         \read_value_mux[5][5] , \read_value_mux[5][4] ,
         \read_value_mux[5][3] , \read_value_mux[5][2] ,
         \read_value_mux[5][1] , \read_value_mux[5][0] ,
         \read_value_mux[4][31] , \read_value_mux[4][30] ,
         \read_value_mux[4][29] , \read_value_mux[4][28] ,
         \read_value_mux[4][27] , \read_value_mux[4][26] ,
         \read_value_mux[4][25] , \read_value_mux[4][24] ,
         \read_value_mux[4][23] , \read_value_mux[4][22] ,
         \read_value_mux[4][21] , \read_value_mux[4][20] ,
         \read_value_mux[4][19] , \read_value_mux[4][18] ,
         \read_value_mux[4][17] , \read_value_mux[4][16] ,
         \read_value_mux[4][15] , \read_value_mux[4][14] ,
         \read_value_mux[4][13] , \read_value_mux[4][12] ,
         \read_value_mux[4][11] , \read_value_mux[4][10] ,
         \read_value_mux[4][9] , \read_value_mux[4][8] ,
         \read_value_mux[4][7] , \read_value_mux[4][6] ,
         \read_value_mux[4][5] , \read_value_mux[4][4] ,
         \read_value_mux[4][3] , \read_value_mux[4][2] ,
         \read_value_mux[4][1] , \read_value_mux[4][0] ,
         \read_value_mux[3][31] , \read_value_mux[3][30] ,
         \read_value_mux[3][29] , \read_value_mux[3][28] ,
         \read_value_mux[3][27] , \read_value_mux[3][26] ,
         \read_value_mux[3][25] , \read_value_mux[3][24] ,
         \read_value_mux[3][23] , \read_value_mux[3][22] ,
         \read_value_mux[3][21] , \read_value_mux[3][20] ,
         \read_value_mux[3][19] , \read_value_mux[3][18] ,
         \read_value_mux[3][17] , \read_value_mux[3][16] ,
         \read_value_mux[3][15] , \read_value_mux[3][14] ,
         \read_value_mux[3][13] , \read_value_mux[3][12] ,
         \read_value_mux[3][11] , \read_value_mux[3][10] ,
         \read_value_mux[3][9] , \read_value_mux[3][8] ,
         \read_value_mux[3][7] , \read_value_mux[3][6] ,
         \read_value_mux[3][5] , \read_value_mux[3][4] ,
         \read_value_mux[3][3] , \read_value_mux[3][2] ,
         \read_value_mux[3][1] , \read_value_mux[3][0] ,
         \read_value_mux[2][31] , \read_value_mux[2][30] ,
         \read_value_mux[2][29] , \read_value_mux[2][28] ,
         \read_value_mux[2][27] , \read_value_mux[2][26] ,
         \read_value_mux[2][25] , \read_value_mux[2][24] ,
         \read_value_mux[2][23] , \read_value_mux[2][22] ,
         \read_value_mux[2][21] , \read_value_mux[2][20] ,
         \read_value_mux[2][19] , \read_value_mux[2][18] ,
         \read_value_mux[2][17] , \read_value_mux[2][16] ,
         \read_value_mux[2][15] , \read_value_mux[2][14] ,
         \read_value_mux[2][13] , \read_value_mux[2][12] ,
         \read_value_mux[2][11] , \read_value_mux[2][10] ,
         \read_value_mux[2][9] , \read_value_mux[2][8] ,
         \read_value_mux[2][7] , \read_value_mux[2][6] ,
         \read_value_mux[2][5] , \read_value_mux[2][4] ,
         \read_value_mux[2][3] , \read_value_mux[2][2] ,
         \read_value_mux[2][1] , \read_value_mux[2][0] ,
         \read_value_mux[1][31] , \read_value_mux[1][30] ,
         \read_value_mux[1][29] , \read_value_mux[1][28] ,
         \read_value_mux[1][27] , \read_value_mux[1][26] ,
         \read_value_mux[1][25] , \read_value_mux[1][24] ,
         \read_value_mux[1][23] , \read_value_mux[1][22] ,
         \read_value_mux[1][21] , \read_value_mux[1][20] ,
         \read_value_mux[1][19] , \read_value_mux[1][18] ,
         \read_value_mux[1][17] , \read_value_mux[1][16] ,
         \read_value_mux[1][15] , \read_value_mux[1][14] ,
         \read_value_mux[1][13] , \read_value_mux[1][12] ,
         \read_value_mux[1][11] , \read_value_mux[1][10] ,
         \read_value_mux[1][9] , \read_value_mux[1][8] ,
         \read_value_mux[1][7] , \read_value_mux[1][6] ,
         \read_value_mux[1][5] , \read_value_mux[1][4] ,
         \read_value_mux[1][3] , \read_value_mux[1][2] ,
         \read_value_mux[1][1] , \read_value_mux[1][0] ,
         \read_value_mux[0][31] , \read_value_mux[0][30] ,
         \read_value_mux[0][29] , \read_value_mux[0][28] ,
         \read_value_mux[0][27] , \read_value_mux[0][26] ,
         \read_value_mux[0][25] , \read_value_mux[0][24] ,
         \read_value_mux[0][23] , \read_value_mux[0][22] ,
         \read_value_mux[0][21] , \read_value_mux[0][20] ,
         \read_value_mux[0][19] , \read_value_mux[0][18] ,
         \read_value_mux[0][17] , \read_value_mux[0][16] ,
         \read_value_mux[0][15] , \read_value_mux[0][14] ,
         \read_value_mux[0][13] , \read_value_mux[0][12] ,
         \read_value_mux[0][11] , \read_value_mux[0][10] ,
         \read_value_mux[0][9] , \read_value_mux[0][8] ,
         \read_value_mux[0][7] , \read_value_mux[0][6] ,
         \read_value_mux[0][5] , \read_value_mux[0][4] ,
         \read_value_mux[0][3] , \read_value_mux[0][2] ,
         \read_value_mux[0][1] , \read_value_mux[0][0] , \words[31]/valid_o ,
         \words[31]/valid_i , \words[31]/data_i[31] , \words[31]/data_i[30] ,
         \words[31]/data_i[29] , \words[31]/data_i[28] ,
         \words[31]/data_i[27] , \words[31]/data_i[26] ,
         \words[31]/data_i[25] , \words[31]/data_i[24] ,
         \words[31]/data_i[23] , \words[31]/data_i[22] ,
         \words[31]/data_i[21] , \words[31]/data_i[20] ,
         \words[31]/data_i[19] , \words[31]/data_i[18] ,
         \words[31]/data_i[17] , \words[31]/data_i[16] ,
         \words[31]/data_i[15] , \words[31]/data_i[14] ,
         \words[31]/data_i[13] , \words[31]/data_i[12] ,
         \words[31]/data_i[11] , \words[31]/data_i[10] , \words[31]/data_i[9] ,
         \words[31]/data_i[8] , \words[31]/data_i[7] , \words[31]/data_i[6] ,
         \words[31]/data_i[5] , \words[31]/data_i[4] , \words[31]/data_i[3] ,
         \words[31]/data_i[2] , \words[31]/data_i[1] , \words[31]/data_i[0] ,
         \words[0]/valid_o , \words[0]/valid_i , \words[0]/data_i[31] ,
         \words[0]/data_i[30] , \words[0]/data_i[29] , \words[0]/data_i[28] ,
         \words[0]/data_i[27] , \words[0]/data_i[26] , \words[0]/data_i[25] ,
         \words[0]/data_i[24] , \words[0]/data_i[23] , \words[0]/data_i[22] ,
         \words[0]/data_i[21] , \words[0]/data_i[20] , \words[0]/data_i[19] ,
         \words[0]/data_i[18] , \words[0]/data_i[17] , \words[0]/data_i[16] ,
         \words[0]/data_i[15] , \words[0]/data_i[14] , \words[0]/data_i[13] ,
         \words[0]/data_i[12] , \words[0]/data_i[11] , \words[0]/data_i[10] ,
         \words[0]/data_i[9] , \words[0]/data_i[8] , \words[0]/data_i[7] ,
         \words[0]/data_i[6] , \words[0]/data_i[5] , \words[0]/data_i[4] ,
         \words[0]/data_i[3] , \words[0]/data_i[2] , \words[0]/data_i[1] ,
         \words[0]/data_i[0] , \words[1]/valid_o , \words[1]/valid_i ,
         \words[1]/data_i[31] , \words[1]/data_i[30] , \words[1]/data_i[29] ,
         \words[1]/data_i[28] , \words[1]/data_i[27] , \words[1]/data_i[26] ,
         \words[1]/data_i[25] , \words[1]/data_i[24] , \words[1]/data_i[23] ,
         \words[1]/data_i[22] , \words[1]/data_i[21] , \words[1]/data_i[20] ,
         \words[1]/data_i[19] , \words[1]/data_i[18] , \words[1]/data_i[17] ,
         \words[1]/data_i[16] , \words[1]/data_i[15] , \words[1]/data_i[14] ,
         \words[1]/data_i[13] , \words[1]/data_i[12] , \words[1]/data_i[11] ,
         \words[1]/data_i[10] , \words[1]/data_i[9] , \words[1]/data_i[8] ,
         \words[1]/data_i[7] , \words[1]/data_i[6] , \words[1]/data_i[5] ,
         \words[1]/data_i[4] , \words[1]/data_i[3] , \words[1]/data_i[2] ,
         \words[1]/data_i[1] , \words[1]/data_i[0] , \words[2]/valid_o ,
         \words[2]/valid_i , \words[2]/data_i[31] , \words[2]/data_i[30] ,
         \words[2]/data_i[29] , \words[2]/data_i[28] , \words[2]/data_i[27] ,
         \words[2]/data_i[26] , \words[2]/data_i[25] , \words[2]/data_i[24] ,
         \words[2]/data_i[23] , \words[2]/data_i[22] , \words[2]/data_i[21] ,
         \words[2]/data_i[20] , \words[2]/data_i[19] , \words[2]/data_i[18] ,
         \words[2]/data_i[17] , \words[2]/data_i[16] , \words[2]/data_i[15] ,
         \words[2]/data_i[14] , \words[2]/data_i[13] , \words[2]/data_i[12] ,
         \words[2]/data_i[11] , \words[2]/data_i[10] , \words[2]/data_i[9] ,
         \words[2]/data_i[8] , \words[2]/data_i[7] , \words[2]/data_i[6] ,
         \words[2]/data_i[5] , \words[2]/data_i[4] , \words[2]/data_i[3] ,
         \words[2]/data_i[2] , \words[2]/data_i[1] , \words[2]/data_i[0] ,
         \words[3]/valid_o , \words[3]/valid_i , \words[3]/data_i[31] ,
         \words[3]/data_i[30] , \words[3]/data_i[29] , \words[3]/data_i[28] ,
         \words[3]/data_i[27] , \words[3]/data_i[26] , \words[3]/data_i[25] ,
         \words[3]/data_i[24] , \words[3]/data_i[23] , \words[3]/data_i[22] ,
         \words[3]/data_i[21] , \words[3]/data_i[20] , \words[3]/data_i[19] ,
         \words[3]/data_i[18] , \words[3]/data_i[17] , \words[3]/data_i[16] ,
         \words[3]/data_i[15] , \words[3]/data_i[14] , \words[3]/data_i[13] ,
         \words[3]/data_i[12] , \words[3]/data_i[11] , \words[3]/data_i[10] ,
         \words[3]/data_i[9] , \words[3]/data_i[8] , \words[3]/data_i[7] ,
         \words[3]/data_i[6] , \words[3]/data_i[5] , \words[3]/data_i[4] ,
         \words[3]/data_i[3] , \words[3]/data_i[2] , \words[3]/data_i[1] ,
         \words[3]/data_i[0] , \words[4]/valid_o , \words[4]/valid_i ,
         \words[4]/data_i[31] , \words[4]/data_i[30] , \words[4]/data_i[29] ,
         \words[4]/data_i[28] , \words[4]/data_i[27] , \words[4]/data_i[26] ,
         \words[4]/data_i[25] , \words[4]/data_i[24] , \words[4]/data_i[23] ,
         \words[4]/data_i[22] , \words[4]/data_i[21] , \words[4]/data_i[20] ,
         \words[4]/data_i[19] , \words[4]/data_i[18] , \words[4]/data_i[17] ,
         \words[4]/data_i[16] , \words[4]/data_i[15] , \words[4]/data_i[14] ,
         \words[4]/data_i[13] , \words[4]/data_i[12] , \words[4]/data_i[11] ,
         \words[4]/data_i[10] , \words[4]/data_i[9] , \words[4]/data_i[8] ,
         \words[4]/data_i[7] , \words[4]/data_i[6] , \words[4]/data_i[5] ,
         \words[4]/data_i[4] , \words[4]/data_i[3] , \words[4]/data_i[2] ,
         \words[4]/data_i[1] , \words[4]/data_i[0] , \words[5]/valid_o ,
         \words[5]/valid_i , \words[5]/data_i[31] , \words[5]/data_i[30] ,
         \words[5]/data_i[29] , \words[5]/data_i[28] , \words[5]/data_i[27] ,
         \words[5]/data_i[26] , \words[5]/data_i[25] , \words[5]/data_i[24] ,
         \words[5]/data_i[23] , \words[5]/data_i[22] , \words[5]/data_i[21] ,
         \words[5]/data_i[20] , \words[5]/data_i[19] , \words[5]/data_i[18] ,
         \words[5]/data_i[17] , \words[5]/data_i[16] , \words[5]/data_i[15] ,
         \words[5]/data_i[14] , \words[5]/data_i[13] , \words[5]/data_i[12] ,
         \words[5]/data_i[11] , \words[5]/data_i[10] , \words[5]/data_i[9] ,
         \words[5]/data_i[8] , \words[5]/data_i[7] , \words[5]/data_i[6] ,
         \words[5]/data_i[5] , \words[5]/data_i[4] , \words[5]/data_i[3] ,
         \words[5]/data_i[2] , \words[5]/data_i[1] , \words[5]/data_i[0] ,
         \words[6]/valid_o , \words[6]/valid_i , \words[6]/data_i[31] ,
         \words[6]/data_i[30] , \words[6]/data_i[29] , \words[6]/data_i[28] ,
         \words[6]/data_i[27] , \words[6]/data_i[26] , \words[6]/data_i[25] ,
         \words[6]/data_i[24] , \words[6]/data_i[23] , \words[6]/data_i[22] ,
         \words[6]/data_i[21] , \words[6]/data_i[20] , \words[6]/data_i[19] ,
         \words[6]/data_i[18] , \words[6]/data_i[17] , \words[6]/data_i[16] ,
         \words[6]/data_i[15] , \words[6]/data_i[14] , \words[6]/data_i[13] ,
         \words[6]/data_i[12] , \words[6]/data_i[11] , \words[6]/data_i[10] ,
         \words[6]/data_i[9] , \words[6]/data_i[8] , \words[6]/data_i[7] ,
         \words[6]/data_i[6] , \words[6]/data_i[5] , \words[6]/data_i[4] ,
         \words[6]/data_i[3] , \words[6]/data_i[2] , \words[6]/data_i[1] ,
         \words[6]/data_i[0] , \words[7]/valid_o , \words[7]/valid_i ,
         \words[7]/data_i[31] , \words[7]/data_i[30] , \words[7]/data_i[29] ,
         \words[7]/data_i[28] , \words[7]/data_i[27] , \words[7]/data_i[26] ,
         \words[7]/data_i[25] , \words[7]/data_i[24] , \words[7]/data_i[23] ,
         \words[7]/data_i[22] , \words[7]/data_i[21] , \words[7]/data_i[20] ,
         \words[7]/data_i[19] , \words[7]/data_i[18] , \words[7]/data_i[17] ,
         \words[7]/data_i[16] , \words[7]/data_i[15] , \words[7]/data_i[14] ,
         \words[7]/data_i[13] , \words[7]/data_i[12] , \words[7]/data_i[11] ,
         \words[7]/data_i[10] , \words[7]/data_i[9] , \words[7]/data_i[8] ,
         \words[7]/data_i[7] , \words[7]/data_i[6] , \words[7]/data_i[5] ,
         \words[7]/data_i[4] , \words[7]/data_i[3] , \words[7]/data_i[2] ,
         \words[7]/data_i[1] , \words[7]/data_i[0] , \words[8]/valid_o ,
         \words[8]/valid_i , \words[8]/data_i[31] , \words[8]/data_i[30] ,
         \words[8]/data_i[29] , \words[8]/data_i[28] , \words[8]/data_i[27] ,
         \words[8]/data_i[26] , \words[8]/data_i[25] , \words[8]/data_i[24] ,
         \words[8]/data_i[23] , \words[8]/data_i[22] , \words[8]/data_i[21] ,
         \words[8]/data_i[20] , \words[8]/data_i[19] , \words[8]/data_i[18] ,
         \words[8]/data_i[17] , \words[8]/data_i[16] , \words[8]/data_i[15] ,
         \words[8]/data_i[14] , \words[8]/data_i[13] , \words[8]/data_i[12] ,
         \words[8]/data_i[11] , \words[8]/data_i[10] , \words[8]/data_i[9] ,
         \words[8]/data_i[8] , \words[8]/data_i[7] , \words[8]/data_i[6] ,
         \words[8]/data_i[5] , \words[8]/data_i[4] , \words[8]/data_i[3] ,
         \words[8]/data_i[2] , \words[8]/data_i[1] , \words[8]/data_i[0] ,
         \words[9]/valid_o , \words[9]/valid_i , \words[9]/data_i[31] ,
         \words[9]/data_i[30] , \words[9]/data_i[29] , \words[9]/data_i[28] ,
         \words[9]/data_i[27] , \words[9]/data_i[26] , \words[9]/data_i[25] ,
         \words[9]/data_i[24] , \words[9]/data_i[23] , \words[9]/data_i[22] ,
         \words[9]/data_i[21] , \words[9]/data_i[20] , \words[9]/data_i[19] ,
         \words[9]/data_i[18] , \words[9]/data_i[17] , \words[9]/data_i[16] ,
         \words[9]/data_i[15] , \words[9]/data_i[14] , \words[9]/data_i[13] ,
         \words[9]/data_i[12] , \words[9]/data_i[11] , \words[9]/data_i[10] ,
         \words[9]/data_i[9] , \words[9]/data_i[8] , \words[9]/data_i[7] ,
         \words[9]/data_i[6] , \words[9]/data_i[5] , \words[9]/data_i[4] ,
         \words[9]/data_i[3] , \words[9]/data_i[2] , \words[9]/data_i[1] ,
         \words[9]/data_i[0] , \words[10]/valid_o , \words[10]/valid_i ,
         \words[10]/data_i[31] , \words[10]/data_i[30] ,
         \words[10]/data_i[29] , \words[10]/data_i[28] ,
         \words[10]/data_i[27] , \words[10]/data_i[26] ,
         \words[10]/data_i[25] , \words[10]/data_i[24] ,
         \words[10]/data_i[23] , \words[10]/data_i[22] ,
         \words[10]/data_i[21] , \words[10]/data_i[20] ,
         \words[10]/data_i[19] , \words[10]/data_i[18] ,
         \words[10]/data_i[17] , \words[10]/data_i[16] ,
         \words[10]/data_i[15] , \words[10]/data_i[14] ,
         \words[10]/data_i[13] , \words[10]/data_i[12] ,
         \words[10]/data_i[11] , \words[10]/data_i[10] , \words[10]/data_i[9] ,
         \words[10]/data_i[8] , \words[10]/data_i[7] , \words[10]/data_i[6] ,
         \words[10]/data_i[5] , \words[10]/data_i[4] , \words[10]/data_i[3] ,
         \words[10]/data_i[2] , \words[10]/data_i[1] , \words[10]/data_i[0] ,
         \words[11]/valid_o , \words[11]/valid_i , \words[11]/data_i[31] ,
         \words[11]/data_i[30] , \words[11]/data_i[29] ,
         \words[11]/data_i[28] , \words[11]/data_i[27] ,
         \words[11]/data_i[26] , \words[11]/data_i[25] ,
         \words[11]/data_i[24] , \words[11]/data_i[23] ,
         \words[11]/data_i[22] , \words[11]/data_i[21] ,
         \words[11]/data_i[20] , \words[11]/data_i[19] ,
         \words[11]/data_i[18] , \words[11]/data_i[17] ,
         \words[11]/data_i[16] , \words[11]/data_i[15] ,
         \words[11]/data_i[14] , \words[11]/data_i[13] ,
         \words[11]/data_i[12] , \words[11]/data_i[11] ,
         \words[11]/data_i[10] , \words[11]/data_i[9] , \words[11]/data_i[8] ,
         \words[11]/data_i[7] , \words[11]/data_i[6] , \words[11]/data_i[5] ,
         \words[11]/data_i[4] , \words[11]/data_i[3] , \words[11]/data_i[2] ,
         \words[11]/data_i[1] , \words[11]/data_i[0] , \words[12]/valid_o ,
         \words[12]/valid_i , \words[12]/data_i[31] , \words[12]/data_i[30] ,
         \words[12]/data_i[29] , \words[12]/data_i[28] ,
         \words[12]/data_i[27] , \words[12]/data_i[26] ,
         \words[12]/data_i[25] , \words[12]/data_i[24] ,
         \words[12]/data_i[23] , \words[12]/data_i[22] ,
         \words[12]/data_i[21] , \words[12]/data_i[20] ,
         \words[12]/data_i[19] , \words[12]/data_i[18] ,
         \words[12]/data_i[17] , \words[12]/data_i[16] ,
         \words[12]/data_i[15] , \words[12]/data_i[14] ,
         \words[12]/data_i[13] , \words[12]/data_i[12] ,
         \words[12]/data_i[11] , \words[12]/data_i[10] , \words[12]/data_i[9] ,
         \words[12]/data_i[8] , \words[12]/data_i[7] , \words[12]/data_i[6] ,
         \words[12]/data_i[5] , \words[12]/data_i[4] , \words[12]/data_i[3] ,
         \words[12]/data_i[2] , \words[12]/data_i[1] , \words[12]/data_i[0] ,
         \words[13]/valid_o , \words[13]/valid_i , \words[13]/data_i[31] ,
         \words[13]/data_i[30] , \words[13]/data_i[29] ,
         \words[13]/data_i[28] , \words[13]/data_i[27] ,
         \words[13]/data_i[26] , \words[13]/data_i[25] ,
         \words[13]/data_i[24] , \words[13]/data_i[23] ,
         \words[13]/data_i[22] , \words[13]/data_i[21] ,
         \words[13]/data_i[20] , \words[13]/data_i[19] ,
         \words[13]/data_i[18] , \words[13]/data_i[17] ,
         \words[13]/data_i[16] , \words[13]/data_i[15] ,
         \words[13]/data_i[14] , \words[13]/data_i[13] ,
         \words[13]/data_i[12] , \words[13]/data_i[11] ,
         \words[13]/data_i[10] , \words[13]/data_i[9] , \words[13]/data_i[8] ,
         \words[13]/data_i[7] , \words[13]/data_i[6] , \words[13]/data_i[5] ,
         \words[13]/data_i[4] , \words[13]/data_i[3] , \words[13]/data_i[2] ,
         \words[13]/data_i[1] , \words[13]/data_i[0] , \words[14]/valid_o ,
         \words[14]/valid_i , \words[14]/data_i[31] , \words[14]/data_i[30] ,
         \words[14]/data_i[29] , \words[14]/data_i[28] ,
         \words[14]/data_i[27] , \words[14]/data_i[26] ,
         \words[14]/data_i[25] , \words[14]/data_i[24] ,
         \words[14]/data_i[23] , \words[14]/data_i[22] ,
         \words[14]/data_i[21] , \words[14]/data_i[20] ,
         \words[14]/data_i[19] , \words[14]/data_i[18] ,
         \words[14]/data_i[17] , \words[14]/data_i[16] ,
         \words[14]/data_i[15] , \words[14]/data_i[14] ,
         \words[14]/data_i[13] , \words[14]/data_i[12] ,
         \words[14]/data_i[11] , \words[14]/data_i[10] , \words[14]/data_i[9] ,
         \words[14]/data_i[8] , \words[14]/data_i[7] , \words[14]/data_i[6] ,
         \words[14]/data_i[5] , \words[14]/data_i[4] , \words[14]/data_i[3] ,
         \words[14]/data_i[2] , \words[14]/data_i[1] , \words[14]/data_i[0] ,
         \words[15]/valid_o , \words[15]/valid_i , \words[15]/data_i[31] ,
         \words[15]/data_i[30] , \words[15]/data_i[29] ,
         \words[15]/data_i[28] , \words[15]/data_i[27] ,
         \words[15]/data_i[26] , \words[15]/data_i[25] ,
         \words[15]/data_i[24] , \words[15]/data_i[23] ,
         \words[15]/data_i[22] , \words[15]/data_i[21] ,
         \words[15]/data_i[20] , \words[15]/data_i[19] ,
         \words[15]/data_i[18] , \words[15]/data_i[17] ,
         \words[15]/data_i[16] , \words[15]/data_i[15] ,
         \words[15]/data_i[14] , \words[15]/data_i[13] ,
         \words[15]/data_i[12] , \words[15]/data_i[11] ,
         \words[15]/data_i[10] , \words[15]/data_i[9] , \words[15]/data_i[8] ,
         \words[15]/data_i[7] , \words[15]/data_i[6] , \words[15]/data_i[5] ,
         \words[15]/data_i[4] , \words[15]/data_i[3] , \words[15]/data_i[2] ,
         \words[15]/data_i[1] , \words[15]/data_i[0] , \words[16]/valid_o ,
         \words[16]/valid_i , \words[16]/data_i[31] , \words[16]/data_i[30] ,
         \words[16]/data_i[29] , \words[16]/data_i[28] ,
         \words[16]/data_i[27] , \words[16]/data_i[26] ,
         \words[16]/data_i[25] , \words[16]/data_i[24] ,
         \words[16]/data_i[23] , \words[16]/data_i[22] ,
         \words[16]/data_i[21] , \words[16]/data_i[20] ,
         \words[16]/data_i[19] , \words[16]/data_i[18] ,
         \words[16]/data_i[17] , \words[16]/data_i[16] ,
         \words[16]/data_i[15] , \words[16]/data_i[14] ,
         \words[16]/data_i[13] , \words[16]/data_i[12] ,
         \words[16]/data_i[11] , \words[16]/data_i[10] , \words[16]/data_i[9] ,
         \words[16]/data_i[8] , \words[16]/data_i[7] , \words[16]/data_i[6] ,
         \words[16]/data_i[5] , \words[16]/data_i[4] , \words[16]/data_i[3] ,
         \words[16]/data_i[2] , \words[16]/data_i[1] , \words[16]/data_i[0] ,
         \words[17]/valid_o , \words[17]/valid_i , \words[17]/data_i[31] ,
         \words[17]/data_i[30] , \words[17]/data_i[29] ,
         \words[17]/data_i[28] , \words[17]/data_i[27] ,
         \words[17]/data_i[26] , \words[17]/data_i[25] ,
         \words[17]/data_i[24] , \words[17]/data_i[23] ,
         \words[17]/data_i[22] , \words[17]/data_i[21] ,
         \words[17]/data_i[20] , \words[17]/data_i[19] ,
         \words[17]/data_i[18] , \words[17]/data_i[17] ,
         \words[17]/data_i[16] , \words[17]/data_i[15] ,
         \words[17]/data_i[14] , \words[17]/data_i[13] ,
         \words[17]/data_i[12] , \words[17]/data_i[11] ,
         \words[17]/data_i[10] , \words[17]/data_i[9] , \words[17]/data_i[8] ,
         \words[17]/data_i[7] , \words[17]/data_i[6] , \words[17]/data_i[5] ,
         \words[17]/data_i[4] , \words[17]/data_i[3] , \words[17]/data_i[2] ,
         \words[17]/data_i[1] , \words[17]/data_i[0] , \words[18]/valid_o ,
         \words[18]/valid_i , \words[18]/data_i[31] , \words[18]/data_i[30] ,
         \words[18]/data_i[29] , \words[18]/data_i[28] ,
         \words[18]/data_i[27] , \words[18]/data_i[26] ,
         \words[18]/data_i[25] , \words[18]/data_i[24] ,
         \words[18]/data_i[23] , \words[18]/data_i[22] ,
         \words[18]/data_i[21] , \words[18]/data_i[20] ,
         \words[18]/data_i[19] , \words[18]/data_i[18] ,
         \words[18]/data_i[17] , \words[18]/data_i[16] ,
         \words[18]/data_i[15] , \words[18]/data_i[14] ,
         \words[18]/data_i[13] , \words[18]/data_i[12] ,
         \words[18]/data_i[11] , \words[18]/data_i[10] , \words[18]/data_i[9] ,
         \words[18]/data_i[8] , \words[18]/data_i[7] , \words[18]/data_i[6] ,
         \words[18]/data_i[5] , \words[18]/data_i[4] , \words[18]/data_i[3] ,
         \words[18]/data_i[2] , \words[18]/data_i[1] , \words[18]/data_i[0] ,
         \words[19]/valid_o , \words[19]/valid_i , \words[19]/data_i[31] ,
         \words[19]/data_i[30] , \words[19]/data_i[29] ,
         \words[19]/data_i[28] , \words[19]/data_i[27] ,
         \words[19]/data_i[26] , \words[19]/data_i[25] ,
         \words[19]/data_i[24] , \words[19]/data_i[23] ,
         \words[19]/data_i[22] , \words[19]/data_i[21] ,
         \words[19]/data_i[20] , \words[19]/data_i[19] ,
         \words[19]/data_i[18] , \words[19]/data_i[17] ,
         \words[19]/data_i[16] , \words[19]/data_i[15] ,
         \words[19]/data_i[14] , \words[19]/data_i[13] ,
         \words[19]/data_i[12] , \words[19]/data_i[11] ,
         \words[19]/data_i[10] , \words[19]/data_i[9] , \words[19]/data_i[8] ,
         \words[19]/data_i[7] , \words[19]/data_i[6] , \words[19]/data_i[5] ,
         \words[19]/data_i[4] , \words[19]/data_i[3] , \words[19]/data_i[2] ,
         \words[19]/data_i[1] , \words[19]/data_i[0] , \words[20]/valid_o ,
         \words[20]/valid_i , \words[20]/data_i[31] , \words[20]/data_i[30] ,
         \words[20]/data_i[29] , \words[20]/data_i[28] ,
         \words[20]/data_i[27] , \words[20]/data_i[26] ,
         \words[20]/data_i[25] , \words[20]/data_i[24] ,
         \words[20]/data_i[23] , \words[20]/data_i[22] ,
         \words[20]/data_i[21] , \words[20]/data_i[20] ,
         \words[20]/data_i[19] , \words[20]/data_i[18] ,
         \words[20]/data_i[17] , \words[20]/data_i[16] ,
         \words[20]/data_i[15] , \words[20]/data_i[14] ,
         \words[20]/data_i[13] , \words[20]/data_i[12] ,
         \words[20]/data_i[11] , \words[20]/data_i[10] , \words[20]/data_i[9] ,
         \words[20]/data_i[8] , \words[20]/data_i[7] , \words[20]/data_i[6] ,
         \words[20]/data_i[5] , \words[20]/data_i[4] , \words[20]/data_i[3] ,
         \words[20]/data_i[2] , \words[20]/data_i[1] , \words[20]/data_i[0] ,
         \words[21]/valid_o , \words[21]/valid_i , \words[21]/data_i[31] ,
         \words[21]/data_i[30] , \words[21]/data_i[29] ,
         \words[21]/data_i[28] , \words[21]/data_i[27] ,
         \words[21]/data_i[26] , \words[21]/data_i[25] ,
         \words[21]/data_i[24] , \words[21]/data_i[23] ,
         \words[21]/data_i[22] , \words[21]/data_i[21] ,
         \words[21]/data_i[20] , \words[21]/data_i[19] ,
         \words[21]/data_i[18] , \words[21]/data_i[17] ,
         \words[21]/data_i[16] , \words[21]/data_i[15] ,
         \words[21]/data_i[14] , \words[21]/data_i[13] ,
         \words[21]/data_i[12] , \words[21]/data_i[11] ,
         \words[21]/data_i[10] , \words[21]/data_i[9] , \words[21]/data_i[8] ,
         \words[21]/data_i[7] , \words[21]/data_i[6] , \words[21]/data_i[5] ,
         \words[21]/data_i[4] , \words[21]/data_i[3] , \words[21]/data_i[2] ,
         \words[21]/data_i[1] , \words[21]/data_i[0] , \words[22]/valid_o ,
         \words[22]/valid_i , \words[22]/data_i[31] , \words[22]/data_i[30] ,
         \words[22]/data_i[29] , \words[22]/data_i[28] ,
         \words[22]/data_i[27] , \words[22]/data_i[26] ,
         \words[22]/data_i[25] , \words[22]/data_i[24] ,
         \words[22]/data_i[23] , \words[22]/data_i[22] ,
         \words[22]/data_i[21] , \words[22]/data_i[20] ,
         \words[22]/data_i[19] , \words[22]/data_i[18] ,
         \words[22]/data_i[17] , \words[22]/data_i[16] ,
         \words[22]/data_i[15] , \words[22]/data_i[14] ,
         \words[22]/data_i[13] , \words[22]/data_i[12] ,
         \words[22]/data_i[11] , \words[22]/data_i[10] , \words[22]/data_i[9] ,
         \words[22]/data_i[8] , \words[22]/data_i[7] , \words[22]/data_i[6] ,
         \words[22]/data_i[5] , \words[22]/data_i[4] , \words[22]/data_i[3] ,
         \words[22]/data_i[2] , \words[22]/data_i[1] , \words[22]/data_i[0] ,
         \words[23]/valid_o , \words[23]/valid_i , \words[23]/data_i[31] ,
         \words[23]/data_i[30] , \words[23]/data_i[29] ,
         \words[23]/data_i[28] , \words[23]/data_i[27] ,
         \words[23]/data_i[26] , \words[23]/data_i[25] ,
         \words[23]/data_i[24] , \words[23]/data_i[23] ,
         \words[23]/data_i[22] , \words[23]/data_i[21] ,
         \words[23]/data_i[20] , \words[23]/data_i[19] ,
         \words[23]/data_i[18] , \words[23]/data_i[17] ,
         \words[23]/data_i[16] , \words[23]/data_i[15] ,
         \words[23]/data_i[14] , \words[23]/data_i[13] ,
         \words[23]/data_i[12] , \words[23]/data_i[11] ,
         \words[23]/data_i[10] , \words[23]/data_i[9] , \words[23]/data_i[8] ,
         \words[23]/data_i[7] , \words[23]/data_i[6] , \words[23]/data_i[5] ,
         \words[23]/data_i[4] , \words[23]/data_i[3] , \words[23]/data_i[2] ,
         \words[23]/data_i[1] , \words[23]/data_i[0] , \words[24]/valid_o ,
         \words[24]/valid_i , \words[24]/data_i[31] , \words[24]/data_i[30] ,
         \words[24]/data_i[29] , \words[24]/data_i[28] ,
         \words[24]/data_i[27] , \words[24]/data_i[26] ,
         \words[24]/data_i[25] , \words[24]/data_i[24] ,
         \words[24]/data_i[23] , \words[24]/data_i[22] ,
         \words[24]/data_i[21] , \words[24]/data_i[20] ,
         \words[24]/data_i[19] , \words[24]/data_i[18] ,
         \words[24]/data_i[17] , \words[24]/data_i[16] ,
         \words[24]/data_i[15] , \words[24]/data_i[14] ,
         \words[24]/data_i[13] , \words[24]/data_i[12] ,
         \words[24]/data_i[11] , \words[24]/data_i[10] , \words[24]/data_i[9] ,
         \words[24]/data_i[8] , \words[24]/data_i[7] , \words[24]/data_i[6] ,
         \words[24]/data_i[5] , \words[24]/data_i[4] , \words[24]/data_i[3] ,
         \words[24]/data_i[2] , \words[24]/data_i[1] , \words[24]/data_i[0] ,
         \words[25]/valid_o , \words[25]/valid_i , \words[25]/data_i[31] ,
         \words[25]/data_i[30] , \words[25]/data_i[29] ,
         \words[25]/data_i[28] , \words[25]/data_i[27] ,
         \words[25]/data_i[26] , \words[25]/data_i[25] ,
         \words[25]/data_i[24] , \words[25]/data_i[23] ,
         \words[25]/data_i[22] , \words[25]/data_i[21] ,
         \words[25]/data_i[20] , \words[25]/data_i[19] ,
         \words[25]/data_i[18] , \words[25]/data_i[17] ,
         \words[25]/data_i[16] , \words[25]/data_i[15] ,
         \words[25]/data_i[14] , \words[25]/data_i[13] ,
         \words[25]/data_i[12] , \words[25]/data_i[11] ,
         \words[25]/data_i[10] , \words[25]/data_i[9] , \words[25]/data_i[8] ,
         \words[25]/data_i[7] , \words[25]/data_i[6] , \words[25]/data_i[5] ,
         \words[25]/data_i[4] , \words[25]/data_i[3] , \words[25]/data_i[2] ,
         \words[25]/data_i[1] , \words[25]/data_i[0] , \words[26]/valid_o ,
         \words[26]/valid_i , \words[26]/data_i[31] , \words[26]/data_i[30] ,
         \words[26]/data_i[29] , \words[26]/data_i[28] ,
         \words[26]/data_i[27] , \words[26]/data_i[26] ,
         \words[26]/data_i[25] , \words[26]/data_i[24] ,
         \words[26]/data_i[23] , \words[26]/data_i[22] ,
         \words[26]/data_i[21] , \words[26]/data_i[20] ,
         \words[26]/data_i[19] , \words[26]/data_i[18] ,
         \words[26]/data_i[17] , \words[26]/data_i[16] ,
         \words[26]/data_i[15] , \words[26]/data_i[14] ,
         \words[26]/data_i[13] , \words[26]/data_i[12] ,
         \words[26]/data_i[11] , \words[26]/data_i[10] , \words[26]/data_i[9] ,
         \words[26]/data_i[8] , \words[26]/data_i[7] , \words[26]/data_i[6] ,
         \words[26]/data_i[5] , \words[26]/data_i[4] , \words[26]/data_i[3] ,
         \words[26]/data_i[2] , \words[26]/data_i[1] , \words[26]/data_i[0] ,
         \words[27]/valid_o , \words[27]/valid_i , \words[27]/data_i[31] ,
         \words[27]/data_i[30] , \words[27]/data_i[29] ,
         \words[27]/data_i[28] , \words[27]/data_i[27] ,
         \words[27]/data_i[26] , \words[27]/data_i[25] ,
         \words[27]/data_i[24] , \words[27]/data_i[23] ,
         \words[27]/data_i[22] , \words[27]/data_i[21] ,
         \words[27]/data_i[20] , \words[27]/data_i[19] ,
         \words[27]/data_i[18] , \words[27]/data_i[17] ,
         \words[27]/data_i[16] , \words[27]/data_i[15] ,
         \words[27]/data_i[14] , \words[27]/data_i[13] ,
         \words[27]/data_i[12] , \words[27]/data_i[11] ,
         \words[27]/data_i[10] , \words[27]/data_i[9] , \words[27]/data_i[8] ,
         \words[27]/data_i[7] , \words[27]/data_i[6] , \words[27]/data_i[5] ,
         \words[27]/data_i[4] , \words[27]/data_i[3] , \words[27]/data_i[2] ,
         \words[27]/data_i[1] , \words[27]/data_i[0] , \words[28]/valid_o ,
         \words[28]/valid_i , \words[28]/data_i[31] , \words[28]/data_i[30] ,
         \words[28]/data_i[29] , \words[28]/data_i[28] ,
         \words[28]/data_i[27] , \words[28]/data_i[26] ,
         \words[28]/data_i[25] , \words[28]/data_i[24] ,
         \words[28]/data_i[23] , \words[28]/data_i[22] ,
         \words[28]/data_i[21] , \words[28]/data_i[20] ,
         \words[28]/data_i[19] , \words[28]/data_i[18] ,
         \words[28]/data_i[17] , \words[28]/data_i[16] ,
         \words[28]/data_i[15] , \words[28]/data_i[14] ,
         \words[28]/data_i[13] , \words[28]/data_i[12] ,
         \words[28]/data_i[11] , \words[28]/data_i[10] , \words[28]/data_i[9] ,
         \words[28]/data_i[8] , \words[28]/data_i[7] , \words[28]/data_i[6] ,
         \words[28]/data_i[5] , \words[28]/data_i[4] , \words[28]/data_i[3] ,
         \words[28]/data_i[2] , \words[28]/data_i[1] , \words[28]/data_i[0] ,
         \words[29]/valid_o , \words[29]/valid_i , \words[29]/data_i[31] ,
         \words[29]/data_i[30] , \words[29]/data_i[29] ,
         \words[29]/data_i[28] , \words[29]/data_i[27] ,
         \words[29]/data_i[26] , \words[29]/data_i[25] ,
         \words[29]/data_i[24] , \words[29]/data_i[23] ,
         \words[29]/data_i[22] , \words[29]/data_i[21] ,
         \words[29]/data_i[20] , \words[29]/data_i[19] ,
         \words[29]/data_i[18] , \words[29]/data_i[17] ,
         \words[29]/data_i[16] , \words[29]/data_i[15] ,
         \words[29]/data_i[14] , \words[29]/data_i[13] ,
         \words[29]/data_i[12] , \words[29]/data_i[11] ,
         \words[29]/data_i[10] , \words[29]/data_i[9] , \words[29]/data_i[8] ,
         \words[29]/data_i[7] , \words[29]/data_i[6] , \words[29]/data_i[5] ,
         \words[29]/data_i[4] , \words[29]/data_i[3] , \words[29]/data_i[2] ,
         \words[29]/data_i[1] , \words[29]/data_i[0] , \words[30]/valid_o ,
         \words[30]/valid_i , \words[30]/data_i[31] , \words[30]/data_i[30] ,
         \words[30]/data_i[29] , \words[30]/data_i[28] ,
         \words[30]/data_i[27] , \words[30]/data_i[26] ,
         \words[30]/data_i[25] , \words[30]/data_i[24] ,
         \words[30]/data_i[23] , \words[30]/data_i[22] ,
         \words[30]/data_i[21] , \words[30]/data_i[20] ,
         \words[30]/data_i[19] , \words[30]/data_i[18] ,
         \words[30]/data_i[17] , \words[30]/data_i[16] ,
         \words[30]/data_i[15] , \words[30]/data_i[14] ,
         \words[30]/data_i[13] , \words[30]/data_i[12] ,
         \words[30]/data_i[11] , \words[30]/data_i[10] , \words[30]/data_i[9] ,
         \words[30]/data_i[8] , \words[30]/data_i[7] , \words[30]/data_i[6] ,
         \words[30]/data_i[5] , \words[30]/data_i[4] , \words[30]/data_i[3] ,
         \words[30]/data_i[2] , \words[30]/data_i[1] , \words[30]/data_i[0] ,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192;

  mux read_mux ( .data_i({\read_value_mux[31][31] , \read_value_mux[31][30] , 
        \read_value_mux[31][29] , \read_value_mux[31][28] , 
        \read_value_mux[31][27] , \read_value_mux[31][26] , 
        \read_value_mux[31][25] , \read_value_mux[31][24] , 
        \read_value_mux[31][23] , \read_value_mux[31][22] , 
        \read_value_mux[31][21] , \read_value_mux[31][20] , 
        \read_value_mux[31][19] , \read_value_mux[31][18] , 
        \read_value_mux[31][17] , \read_value_mux[31][16] , 
        \read_value_mux[31][15] , \read_value_mux[31][14] , 
        \read_value_mux[31][13] , \read_value_mux[31][12] , 
        \read_value_mux[31][11] , \read_value_mux[31][10] , 
        \read_value_mux[31][9] , \read_value_mux[31][8] , 
        \read_value_mux[31][7] , \read_value_mux[31][6] , 
        \read_value_mux[31][5] , \read_value_mux[31][4] , 
        \read_value_mux[31][3] , \read_value_mux[31][2] , 
        \read_value_mux[31][1] , \read_value_mux[31][0] , 
        \read_value_mux[30][31] , \read_value_mux[30][30] , 
        \read_value_mux[30][29] , \read_value_mux[30][28] , 
        \read_value_mux[30][27] , \read_value_mux[30][26] , 
        \read_value_mux[30][25] , \read_value_mux[30][24] , 
        \read_value_mux[30][23] , \read_value_mux[30][22] , 
        \read_value_mux[30][21] , \read_value_mux[30][20] , 
        \read_value_mux[30][19] , \read_value_mux[30][18] , 
        \read_value_mux[30][17] , \read_value_mux[30][16] , 
        \read_value_mux[30][15] , \read_value_mux[30][14] , 
        \read_value_mux[30][13] , \read_value_mux[30][12] , 
        \read_value_mux[30][11] , \read_value_mux[30][10] , 
        \read_value_mux[30][9] , \read_value_mux[30][8] , 
        \read_value_mux[30][7] , \read_value_mux[30][6] , 
        \read_value_mux[30][5] , \read_value_mux[30][4] , 
        \read_value_mux[30][3] , \read_value_mux[30][2] , 
        \read_value_mux[30][1] , \read_value_mux[30][0] , 
        \read_value_mux[29][31] , \read_value_mux[29][30] , 
        \read_value_mux[29][29] , \read_value_mux[29][28] , 
        \read_value_mux[29][27] , \read_value_mux[29][26] , 
        \read_value_mux[29][25] , \read_value_mux[29][24] , 
        \read_value_mux[29][23] , \read_value_mux[29][22] , 
        \read_value_mux[29][21] , \read_value_mux[29][20] , 
        \read_value_mux[29][19] , \read_value_mux[29][18] , 
        \read_value_mux[29][17] , \read_value_mux[29][16] , 
        \read_value_mux[29][15] , \read_value_mux[29][14] , 
        \read_value_mux[29][13] , \read_value_mux[29][12] , 
        \read_value_mux[29][11] , \read_value_mux[29][10] , 
        \read_value_mux[29][9] , \read_value_mux[29][8] , 
        \read_value_mux[29][7] , \read_value_mux[29][6] , 
        \read_value_mux[29][5] , \read_value_mux[29][4] , 
        \read_value_mux[29][3] , \read_value_mux[29][2] , 
        \read_value_mux[29][1] , \read_value_mux[29][0] , 
        \read_value_mux[28][31] , \read_value_mux[28][30] , 
        \read_value_mux[28][29] , \read_value_mux[28][28] , 
        \read_value_mux[28][27] , \read_value_mux[28][26] , 
        \read_value_mux[28][25] , \read_value_mux[28][24] , 
        \read_value_mux[28][23] , \read_value_mux[28][22] , 
        \read_value_mux[28][21] , \read_value_mux[28][20] , 
        \read_value_mux[28][19] , \read_value_mux[28][18] , 
        \read_value_mux[28][17] , \read_value_mux[28][16] , 
        \read_value_mux[28][15] , \read_value_mux[28][14] , 
        \read_value_mux[28][13] , \read_value_mux[28][12] , 
        \read_value_mux[28][11] , \read_value_mux[28][10] , 
        \read_value_mux[28][9] , \read_value_mux[28][8] , 
        \read_value_mux[28][7] , \read_value_mux[28][6] , 
        \read_value_mux[28][5] , \read_value_mux[28][4] , 
        \read_value_mux[28][3] , \read_value_mux[28][2] , 
        \read_value_mux[28][1] , \read_value_mux[28][0] , 
        \read_value_mux[27][31] , \read_value_mux[27][30] , 
        \read_value_mux[27][29] , \read_value_mux[27][28] , 
        \read_value_mux[27][27] , \read_value_mux[27][26] , 
        \read_value_mux[27][25] , \read_value_mux[27][24] , 
        \read_value_mux[27][23] , \read_value_mux[27][22] , 
        \read_value_mux[27][21] , \read_value_mux[27][20] , 
        \read_value_mux[27][19] , \read_value_mux[27][18] , 
        \read_value_mux[27][17] , \read_value_mux[27][16] , 
        \read_value_mux[27][15] , \read_value_mux[27][14] , 
        \read_value_mux[27][13] , \read_value_mux[27][12] , 
        \read_value_mux[27][11] , \read_value_mux[27][10] , 
        \read_value_mux[27][9] , \read_value_mux[27][8] , 
        \read_value_mux[27][7] , \read_value_mux[27][6] , 
        \read_value_mux[27][5] , \read_value_mux[27][4] , 
        \read_value_mux[27][3] , \read_value_mux[27][2] , 
        \read_value_mux[27][1] , \read_value_mux[27][0] , 
        \read_value_mux[26][31] , \read_value_mux[26][30] , 
        \read_value_mux[26][29] , \read_value_mux[26][28] , 
        \read_value_mux[26][27] , \read_value_mux[26][26] , 
        \read_value_mux[26][25] , \read_value_mux[26][24] , 
        \read_value_mux[26][23] , \read_value_mux[26][22] , 
        \read_value_mux[26][21] , \read_value_mux[26][20] , 
        \read_value_mux[26][19] , \read_value_mux[26][18] , 
        \read_value_mux[26][17] , \read_value_mux[26][16] , 
        \read_value_mux[26][15] , \read_value_mux[26][14] , 
        \read_value_mux[26][13] , \read_value_mux[26][12] , 
        \read_value_mux[26][11] , \read_value_mux[26][10] , 
        \read_value_mux[26][9] , \read_value_mux[26][8] , 
        \read_value_mux[26][7] , \read_value_mux[26][6] , 
        \read_value_mux[26][5] , \read_value_mux[26][4] , 
        \read_value_mux[26][3] , \read_value_mux[26][2] , 
        \read_value_mux[26][1] , \read_value_mux[26][0] , 
        \read_value_mux[25][31] , \read_value_mux[25][30] , 
        \read_value_mux[25][29] , \read_value_mux[25][28] , 
        \read_value_mux[25][27] , \read_value_mux[25][26] , 
        \read_value_mux[25][25] , \read_value_mux[25][24] , 
        \read_value_mux[25][23] , \read_value_mux[25][22] , 
        \read_value_mux[25][21] , \read_value_mux[25][20] , 
        \read_value_mux[25][19] , \read_value_mux[25][18] , 
        \read_value_mux[25][17] , \read_value_mux[25][16] , 
        \read_value_mux[25][15] , \read_value_mux[25][14] , 
        \read_value_mux[25][13] , \read_value_mux[25][12] , 
        \read_value_mux[25][11] , \read_value_mux[25][10] , 
        \read_value_mux[25][9] , \read_value_mux[25][8] , 
        \read_value_mux[25][7] , \read_value_mux[25][6] , 
        \read_value_mux[25][5] , \read_value_mux[25][4] , 
        \read_value_mux[25][3] , \read_value_mux[25][2] , 
        \read_value_mux[25][1] , \read_value_mux[25][0] , 
        \read_value_mux[24][31] , \read_value_mux[24][30] , 
        \read_value_mux[24][29] , \read_value_mux[24][28] , 
        \read_value_mux[24][27] , \read_value_mux[24][26] , 
        \read_value_mux[24][25] , \read_value_mux[24][24] , 
        \read_value_mux[24][23] , \read_value_mux[24][22] , 
        \read_value_mux[24][21] , \read_value_mux[24][20] , 
        \read_value_mux[24][19] , \read_value_mux[24][18] , 
        \read_value_mux[24][17] , \read_value_mux[24][16] , 
        \read_value_mux[24][15] , \read_value_mux[24][14] , 
        \read_value_mux[24][13] , \read_value_mux[24][12] , 
        \read_value_mux[24][11] , \read_value_mux[24][10] , 
        \read_value_mux[24][9] , \read_value_mux[24][8] , 
        \read_value_mux[24][7] , \read_value_mux[24][6] , 
        \read_value_mux[24][5] , \read_value_mux[24][4] , 
        \read_value_mux[24][3] , \read_value_mux[24][2] , 
        \read_value_mux[24][1] , \read_value_mux[24][0] , 
        \read_value_mux[23][31] , \read_value_mux[23][30] , 
        \read_value_mux[23][29] , \read_value_mux[23][28] , 
        \read_value_mux[23][27] , \read_value_mux[23][26] , 
        \read_value_mux[23][25] , \read_value_mux[23][24] , 
        \read_value_mux[23][23] , \read_value_mux[23][22] , 
        \read_value_mux[23][21] , \read_value_mux[23][20] , 
        \read_value_mux[23][19] , \read_value_mux[23][18] , 
        \read_value_mux[23][17] , \read_value_mux[23][16] , 
        \read_value_mux[23][15] , \read_value_mux[23][14] , 
        \read_value_mux[23][13] , \read_value_mux[23][12] , 
        \read_value_mux[23][11] , \read_value_mux[23][10] , 
        \read_value_mux[23][9] , \read_value_mux[23][8] , 
        \read_value_mux[23][7] , \read_value_mux[23][6] , 
        \read_value_mux[23][5] , \read_value_mux[23][4] , 
        \read_value_mux[23][3] , \read_value_mux[23][2] , 
        \read_value_mux[23][1] , \read_value_mux[23][0] , 
        \read_value_mux[22][31] , \read_value_mux[22][30] , 
        \read_value_mux[22][29] , \read_value_mux[22][28] , 
        \read_value_mux[22][27] , \read_value_mux[22][26] , 
        \read_value_mux[22][25] , \read_value_mux[22][24] , 
        \read_value_mux[22][23] , \read_value_mux[22][22] , 
        \read_value_mux[22][21] , \read_value_mux[22][20] , 
        \read_value_mux[22][19] , \read_value_mux[22][18] , 
        \read_value_mux[22][17] , \read_value_mux[22][16] , 
        \read_value_mux[22][15] , \read_value_mux[22][14] , 
        \read_value_mux[22][13] , \read_value_mux[22][12] , 
        \read_value_mux[22][11] , \read_value_mux[22][10] , 
        \read_value_mux[22][9] , \read_value_mux[22][8] , 
        \read_value_mux[22][7] , \read_value_mux[22][6] , 
        \read_value_mux[22][5] , \read_value_mux[22][4] , 
        \read_value_mux[22][3] , \read_value_mux[22][2] , 
        \read_value_mux[22][1] , \read_value_mux[22][0] , 
        \read_value_mux[21][31] , \read_value_mux[21][30] , 
        \read_value_mux[21][29] , \read_value_mux[21][28] , 
        \read_value_mux[21][27] , \read_value_mux[21][26] , 
        \read_value_mux[21][25] , \read_value_mux[21][24] , 
        \read_value_mux[21][23] , \read_value_mux[21][22] , 
        \read_value_mux[21][21] , \read_value_mux[21][20] , 
        \read_value_mux[21][19] , \read_value_mux[21][18] , 
        \read_value_mux[21][17] , \read_value_mux[21][16] , 
        \read_value_mux[21][15] , \read_value_mux[21][14] , 
        \read_value_mux[21][13] , \read_value_mux[21][12] , 
        \read_value_mux[21][11] , \read_value_mux[21][10] , 
        \read_value_mux[21][9] , \read_value_mux[21][8] , 
        \read_value_mux[21][7] , \read_value_mux[21][6] , 
        \read_value_mux[21][5] , \read_value_mux[21][4] , 
        \read_value_mux[21][3] , \read_value_mux[21][2] , 
        \read_value_mux[21][1] , \read_value_mux[21][0] , 
        \read_value_mux[20][31] , \read_value_mux[20][30] , 
        \read_value_mux[20][29] , \read_value_mux[20][28] , 
        \read_value_mux[20][27] , \read_value_mux[20][26] , 
        \read_value_mux[20][25] , \read_value_mux[20][24] , 
        \read_value_mux[20][23] , \read_value_mux[20][22] , 
        \read_value_mux[20][21] , \read_value_mux[20][20] , 
        \read_value_mux[20][19] , \read_value_mux[20][18] , 
        \read_value_mux[20][17] , \read_value_mux[20][16] , 
        \read_value_mux[20][15] , \read_value_mux[20][14] , 
        \read_value_mux[20][13] , \read_value_mux[20][12] , 
        \read_value_mux[20][11] , \read_value_mux[20][10] , 
        \read_value_mux[20][9] , \read_value_mux[20][8] , 
        \read_value_mux[20][7] , \read_value_mux[20][6] , 
        \read_value_mux[20][5] , \read_value_mux[20][4] , 
        \read_value_mux[20][3] , \read_value_mux[20][2] , 
        \read_value_mux[20][1] , \read_value_mux[20][0] , 
        \read_value_mux[19][31] , \read_value_mux[19][30] , 
        \read_value_mux[19][29] , \read_value_mux[19][28] , 
        \read_value_mux[19][27] , \read_value_mux[19][26] , 
        \read_value_mux[19][25] , \read_value_mux[19][24] , 
        \read_value_mux[19][23] , \read_value_mux[19][22] , 
        \read_value_mux[19][21] , \read_value_mux[19][20] , 
        \read_value_mux[19][19] , \read_value_mux[19][18] , 
        \read_value_mux[19][17] , \read_value_mux[19][16] , 
        \read_value_mux[19][15] , \read_value_mux[19][14] , 
        \read_value_mux[19][13] , \read_value_mux[19][12] , 
        \read_value_mux[19][11] , \read_value_mux[19][10] , 
        \read_value_mux[19][9] , \read_value_mux[19][8] , 
        \read_value_mux[19][7] , \read_value_mux[19][6] , 
        \read_value_mux[19][5] , \read_value_mux[19][4] , 
        \read_value_mux[19][3] , \read_value_mux[19][2] , 
        \read_value_mux[19][1] , \read_value_mux[19][0] , 
        \read_value_mux[18][31] , \read_value_mux[18][30] , 
        \read_value_mux[18][29] , \read_value_mux[18][28] , 
        \read_value_mux[18][27] , \read_value_mux[18][26] , 
        \read_value_mux[18][25] , \read_value_mux[18][24] , 
        \read_value_mux[18][23] , \read_value_mux[18][22] , 
        \read_value_mux[18][21] , \read_value_mux[18][20] , 
        \read_value_mux[18][19] , \read_value_mux[18][18] , 
        \read_value_mux[18][17] , \read_value_mux[18][16] , 
        \read_value_mux[18][15] , \read_value_mux[18][14] , 
        \read_value_mux[18][13] , \read_value_mux[18][12] , 
        \read_value_mux[18][11] , \read_value_mux[18][10] , 
        \read_value_mux[18][9] , \read_value_mux[18][8] , 
        \read_value_mux[18][7] , \read_value_mux[18][6] , 
        \read_value_mux[18][5] , \read_value_mux[18][4] , 
        \read_value_mux[18][3] , \read_value_mux[18][2] , 
        \read_value_mux[18][1] , \read_value_mux[18][0] , 
        \read_value_mux[17][31] , \read_value_mux[17][30] , 
        \read_value_mux[17][29] , \read_value_mux[17][28] , 
        \read_value_mux[17][27] , \read_value_mux[17][26] , 
        \read_value_mux[17][25] , \read_value_mux[17][24] , 
        \read_value_mux[17][23] , \read_value_mux[17][22] , 
        \read_value_mux[17][21] , \read_value_mux[17][20] , 
        \read_value_mux[17][19] , \read_value_mux[17][18] , 
        \read_value_mux[17][17] , \read_value_mux[17][16] , 
        \read_value_mux[17][15] , \read_value_mux[17][14] , 
        \read_value_mux[17][13] , \read_value_mux[17][12] , 
        \read_value_mux[17][11] , \read_value_mux[17][10] , 
        \read_value_mux[17][9] , \read_value_mux[17][8] , 
        \read_value_mux[17][7] , \read_value_mux[17][6] , 
        \read_value_mux[17][5] , \read_value_mux[17][4] , 
        \read_value_mux[17][3] , \read_value_mux[17][2] , 
        \read_value_mux[17][1] , \read_value_mux[17][0] , 
        \read_value_mux[16][31] , \read_value_mux[16][30] , 
        \read_value_mux[16][29] , \read_value_mux[16][28] , 
        \read_value_mux[16][27] , \read_value_mux[16][26] , 
        \read_value_mux[16][25] , \read_value_mux[16][24] , 
        \read_value_mux[16][23] , \read_value_mux[16][22] , 
        \read_value_mux[16][21] , \read_value_mux[16][20] , 
        \read_value_mux[16][19] , \read_value_mux[16][18] , 
        \read_value_mux[16][17] , \read_value_mux[16][16] , 
        \read_value_mux[16][15] , \read_value_mux[16][14] , 
        \read_value_mux[16][13] , \read_value_mux[16][12] , 
        \read_value_mux[16][11] , \read_value_mux[16][10] , 
        \read_value_mux[16][9] , \read_value_mux[16][8] , 
        \read_value_mux[16][7] , \read_value_mux[16][6] , 
        \read_value_mux[16][5] , \read_value_mux[16][4] , 
        \read_value_mux[16][3] , \read_value_mux[16][2] , 
        \read_value_mux[16][1] , \read_value_mux[16][0] , 
        \read_value_mux[15][31] , \read_value_mux[15][30] , 
        \read_value_mux[15][29] , \read_value_mux[15][28] , 
        \read_value_mux[15][27] , \read_value_mux[15][26] , 
        \read_value_mux[15][25] , \read_value_mux[15][24] , 
        \read_value_mux[15][23] , \read_value_mux[15][22] , 
        \read_value_mux[15][21] , \read_value_mux[15][20] , 
        \read_value_mux[15][19] , \read_value_mux[15][18] , 
        \read_value_mux[15][17] , \read_value_mux[15][16] , 
        \read_value_mux[15][15] , \read_value_mux[15][14] , 
        \read_value_mux[15][13] , \read_value_mux[15][12] , 
        \read_value_mux[15][11] , \read_value_mux[15][10] , 
        \read_value_mux[15][9] , \read_value_mux[15][8] , 
        \read_value_mux[15][7] , \read_value_mux[15][6] , 
        \read_value_mux[15][5] , \read_value_mux[15][4] , 
        \read_value_mux[15][3] , \read_value_mux[15][2] , 
        \read_value_mux[15][1] , \read_value_mux[15][0] , 
        \read_value_mux[14][31] , \read_value_mux[14][30] , 
        \read_value_mux[14][29] , \read_value_mux[14][28] , 
        \read_value_mux[14][27] , \read_value_mux[14][26] , 
        \read_value_mux[14][25] , \read_value_mux[14][24] , 
        \read_value_mux[14][23] , \read_value_mux[14][22] , 
        \read_value_mux[14][21] , \read_value_mux[14][20] , 
        \read_value_mux[14][19] , \read_value_mux[14][18] , 
        \read_value_mux[14][17] , \read_value_mux[14][16] , 
        \read_value_mux[14][15] , \read_value_mux[14][14] , 
        \read_value_mux[14][13] , \read_value_mux[14][12] , 
        \read_value_mux[14][11] , \read_value_mux[14][10] , 
        \read_value_mux[14][9] , \read_value_mux[14][8] , 
        \read_value_mux[14][7] , \read_value_mux[14][6] , 
        \read_value_mux[14][5] , \read_value_mux[14][4] , 
        \read_value_mux[14][3] , \read_value_mux[14][2] , 
        \read_value_mux[14][1] , \read_value_mux[14][0] , 
        \read_value_mux[13][31] , \read_value_mux[13][30] , 
        \read_value_mux[13][29] , \read_value_mux[13][28] , 
        \read_value_mux[13][27] , \read_value_mux[13][26] , 
        \read_value_mux[13][25] , \read_value_mux[13][24] , 
        \read_value_mux[13][23] , \read_value_mux[13][22] , 
        \read_value_mux[13][21] , \read_value_mux[13][20] , 
        \read_value_mux[13][19] , \read_value_mux[13][18] , 
        \read_value_mux[13][17] , \read_value_mux[13][16] , 
        \read_value_mux[13][15] , \read_value_mux[13][14] , 
        \read_value_mux[13][13] , \read_value_mux[13][12] , 
        \read_value_mux[13][11] , \read_value_mux[13][10] , 
        \read_value_mux[13][9] , \read_value_mux[13][8] , 
        \read_value_mux[13][7] , \read_value_mux[13][6] , 
        \read_value_mux[13][5] , \read_value_mux[13][4] , 
        \read_value_mux[13][3] , \read_value_mux[13][2] , 
        \read_value_mux[13][1] , \read_value_mux[13][0] , 
        \read_value_mux[12][31] , \read_value_mux[12][30] , 
        \read_value_mux[12][29] , \read_value_mux[12][28] , 
        \read_value_mux[12][27] , \read_value_mux[12][26] , 
        \read_value_mux[12][25] , \read_value_mux[12][24] , 
        \read_value_mux[12][23] , \read_value_mux[12][22] , 
        \read_value_mux[12][21] , \read_value_mux[12][20] , 
        \read_value_mux[12][19] , \read_value_mux[12][18] , 
        \read_value_mux[12][17] , \read_value_mux[12][16] , 
        \read_value_mux[12][15] , \read_value_mux[12][14] , 
        \read_value_mux[12][13] , \read_value_mux[12][12] , 
        \read_value_mux[12][11] , \read_value_mux[12][10] , 
        \read_value_mux[12][9] , \read_value_mux[12][8] , 
        \read_value_mux[12][7] , \read_value_mux[12][6] , 
        \read_value_mux[12][5] , \read_value_mux[12][4] , 
        \read_value_mux[12][3] , \read_value_mux[12][2] , 
        \read_value_mux[12][1] , \read_value_mux[12][0] , 
        \read_value_mux[11][31] , \read_value_mux[11][30] , 
        \read_value_mux[11][29] , \read_value_mux[11][28] , 
        \read_value_mux[11][27] , \read_value_mux[11][26] , 
        \read_value_mux[11][25] , \read_value_mux[11][24] , 
        \read_value_mux[11][23] , \read_value_mux[11][22] , 
        \read_value_mux[11][21] , \read_value_mux[11][20] , 
        \read_value_mux[11][19] , \read_value_mux[11][18] , 
        \read_value_mux[11][17] , \read_value_mux[11][16] , 
        \read_value_mux[11][15] , \read_value_mux[11][14] , 
        \read_value_mux[11][13] , \read_value_mux[11][12] , 
        \read_value_mux[11][11] , \read_value_mux[11][10] , 
        \read_value_mux[11][9] , \read_value_mux[11][8] , 
        \read_value_mux[11][7] , \read_value_mux[11][6] , 
        \read_value_mux[11][5] , \read_value_mux[11][4] , 
        \read_value_mux[11][3] , \read_value_mux[11][2] , 
        \read_value_mux[11][1] , \read_value_mux[11][0] , 
        \read_value_mux[10][31] , \read_value_mux[10][30] , 
        \read_value_mux[10][29] , \read_value_mux[10][28] , 
        \read_value_mux[10][27] , \read_value_mux[10][26] , 
        \read_value_mux[10][25] , \read_value_mux[10][24] , 
        \read_value_mux[10][23] , \read_value_mux[10][22] , 
        \read_value_mux[10][21] , \read_value_mux[10][20] , 
        \read_value_mux[10][19] , \read_value_mux[10][18] , 
        \read_value_mux[10][17] , \read_value_mux[10][16] , 
        \read_value_mux[10][15] , \read_value_mux[10][14] , 
        \read_value_mux[10][13] , \read_value_mux[10][12] , 
        \read_value_mux[10][11] , \read_value_mux[10][10] , 
        \read_value_mux[10][9] , \read_value_mux[10][8] , 
        \read_value_mux[10][7] , \read_value_mux[10][6] , 
        \read_value_mux[10][5] , \read_value_mux[10][4] , 
        \read_value_mux[10][3] , \read_value_mux[10][2] , 
        \read_value_mux[10][1] , \read_value_mux[10][0] , 
        \read_value_mux[9][31] , \read_value_mux[9][30] , 
        \read_value_mux[9][29] , \read_value_mux[9][28] , 
        \read_value_mux[9][27] , \read_value_mux[9][26] , 
        \read_value_mux[9][25] , \read_value_mux[9][24] , 
        \read_value_mux[9][23] , \read_value_mux[9][22] , 
        \read_value_mux[9][21] , \read_value_mux[9][20] , 
        \read_value_mux[9][19] , \read_value_mux[9][18] , 
        \read_value_mux[9][17] , \read_value_mux[9][16] , 
        \read_value_mux[9][15] , \read_value_mux[9][14] , 
        \read_value_mux[9][13] , \read_value_mux[9][12] , 
        \read_value_mux[9][11] , \read_value_mux[9][10] , 
        \read_value_mux[9][9] , \read_value_mux[9][8] , \read_value_mux[9][7] , 
        \read_value_mux[9][6] , \read_value_mux[9][5] , \read_value_mux[9][4] , 
        \read_value_mux[9][3] , \read_value_mux[9][2] , \read_value_mux[9][1] , 
        \read_value_mux[9][0] , \read_value_mux[8][31] , 
        \read_value_mux[8][30] , \read_value_mux[8][29] , 
        \read_value_mux[8][28] , \read_value_mux[8][27] , 
        \read_value_mux[8][26] , \read_value_mux[8][25] , 
        \read_value_mux[8][24] , \read_value_mux[8][23] , 
        \read_value_mux[8][22] , \read_value_mux[8][21] , 
        \read_value_mux[8][20] , \read_value_mux[8][19] , 
        \read_value_mux[8][18] , \read_value_mux[8][17] , 
        \read_value_mux[8][16] , \read_value_mux[8][15] , 
        \read_value_mux[8][14] , \read_value_mux[8][13] , 
        \read_value_mux[8][12] , \read_value_mux[8][11] , 
        \read_value_mux[8][10] , \read_value_mux[8][9] , 
        \read_value_mux[8][8] , \read_value_mux[8][7] , \read_value_mux[8][6] , 
        \read_value_mux[8][5] , \read_value_mux[8][4] , \read_value_mux[8][3] , 
        \read_value_mux[8][2] , \read_value_mux[8][1] , \read_value_mux[8][0] , 
        \read_value_mux[7][31] , \read_value_mux[7][30] , 
        \read_value_mux[7][29] , \read_value_mux[7][28] , 
        \read_value_mux[7][27] , \read_value_mux[7][26] , 
        \read_value_mux[7][25] , \read_value_mux[7][24] , 
        \read_value_mux[7][23] , \read_value_mux[7][22] , 
        \read_value_mux[7][21] , \read_value_mux[7][20] , 
        \read_value_mux[7][19] , \read_value_mux[7][18] , 
        \read_value_mux[7][17] , \read_value_mux[7][16] , 
        \read_value_mux[7][15] , \read_value_mux[7][14] , 
        \read_value_mux[7][13] , \read_value_mux[7][12] , 
        \read_value_mux[7][11] , \read_value_mux[7][10] , 
        \read_value_mux[7][9] , \read_value_mux[7][8] , \read_value_mux[7][7] , 
        \read_value_mux[7][6] , \read_value_mux[7][5] , \read_value_mux[7][4] , 
        \read_value_mux[7][3] , \read_value_mux[7][2] , \read_value_mux[7][1] , 
        \read_value_mux[7][0] , \read_value_mux[6][31] , 
        \read_value_mux[6][30] , \read_value_mux[6][29] , 
        \read_value_mux[6][28] , \read_value_mux[6][27] , 
        \read_value_mux[6][26] , \read_value_mux[6][25] , 
        \read_value_mux[6][24] , \read_value_mux[6][23] , 
        \read_value_mux[6][22] , \read_value_mux[6][21] , 
        \read_value_mux[6][20] , \read_value_mux[6][19] , 
        \read_value_mux[6][18] , \read_value_mux[6][17] , 
        \read_value_mux[6][16] , \read_value_mux[6][15] , 
        \read_value_mux[6][14] , \read_value_mux[6][13] , 
        \read_value_mux[6][12] , \read_value_mux[6][11] , 
        \read_value_mux[6][10] , \read_value_mux[6][9] , 
        \read_value_mux[6][8] , \read_value_mux[6][7] , \read_value_mux[6][6] , 
        \read_value_mux[6][5] , \read_value_mux[6][4] , \read_value_mux[6][3] , 
        \read_value_mux[6][2] , \read_value_mux[6][1] , \read_value_mux[6][0] , 
        \read_value_mux[5][31] , \read_value_mux[5][30] , 
        \read_value_mux[5][29] , \read_value_mux[5][28] , 
        \read_value_mux[5][27] , \read_value_mux[5][26] , 
        \read_value_mux[5][25] , \read_value_mux[5][24] , 
        \read_value_mux[5][23] , \read_value_mux[5][22] , 
        \read_value_mux[5][21] , \read_value_mux[5][20] , 
        \read_value_mux[5][19] , \read_value_mux[5][18] , 
        \read_value_mux[5][17] , \read_value_mux[5][16] , 
        \read_value_mux[5][15] , \read_value_mux[5][14] , 
        \read_value_mux[5][13] , \read_value_mux[5][12] , 
        \read_value_mux[5][11] , \read_value_mux[5][10] , 
        \read_value_mux[5][9] , \read_value_mux[5][8] , \read_value_mux[5][7] , 
        \read_value_mux[5][6] , \read_value_mux[5][5] , \read_value_mux[5][4] , 
        \read_value_mux[5][3] , \read_value_mux[5][2] , \read_value_mux[5][1] , 
        \read_value_mux[5][0] , \read_value_mux[4][31] , 
        \read_value_mux[4][30] , \read_value_mux[4][29] , 
        \read_value_mux[4][28] , \read_value_mux[4][27] , 
        \read_value_mux[4][26] , \read_value_mux[4][25] , 
        \read_value_mux[4][24] , \read_value_mux[4][23] , 
        \read_value_mux[4][22] , \read_value_mux[4][21] , 
        \read_value_mux[4][20] , \read_value_mux[4][19] , 
        \read_value_mux[4][18] , \read_value_mux[4][17] , 
        \read_value_mux[4][16] , \read_value_mux[4][15] , 
        \read_value_mux[4][14] , \read_value_mux[4][13] , 
        \read_value_mux[4][12] , \read_value_mux[4][11] , 
        \read_value_mux[4][10] , \read_value_mux[4][9] , 
        \read_value_mux[4][8] , \read_value_mux[4][7] , \read_value_mux[4][6] , 
        \read_value_mux[4][5] , \read_value_mux[4][4] , \read_value_mux[4][3] , 
        \read_value_mux[4][2] , \read_value_mux[4][1] , \read_value_mux[4][0] , 
        \read_value_mux[3][31] , \read_value_mux[3][30] , 
        \read_value_mux[3][29] , \read_value_mux[3][28] , 
        \read_value_mux[3][27] , \read_value_mux[3][26] , 
        \read_value_mux[3][25] , \read_value_mux[3][24] , 
        \read_value_mux[3][23] , \read_value_mux[3][22] , 
        \read_value_mux[3][21] , \read_value_mux[3][20] , 
        \read_value_mux[3][19] , \read_value_mux[3][18] , 
        \read_value_mux[3][17] , \read_value_mux[3][16] , 
        \read_value_mux[3][15] , \read_value_mux[3][14] , 
        \read_value_mux[3][13] , \read_value_mux[3][12] , 
        \read_value_mux[3][11] , \read_value_mux[3][10] , 
        \read_value_mux[3][9] , \read_value_mux[3][8] , \read_value_mux[3][7] , 
        \read_value_mux[3][6] , \read_value_mux[3][5] , \read_value_mux[3][4] , 
        \read_value_mux[3][3] , \read_value_mux[3][2] , \read_value_mux[3][1] , 
        \read_value_mux[3][0] , \read_value_mux[2][31] , 
        \read_value_mux[2][30] , \read_value_mux[2][29] , 
        \read_value_mux[2][28] , \read_value_mux[2][27] , 
        \read_value_mux[2][26] , \read_value_mux[2][25] , 
        \read_value_mux[2][24] , \read_value_mux[2][23] , 
        \read_value_mux[2][22] , \read_value_mux[2][21] , 
        \read_value_mux[2][20] , \read_value_mux[2][19] , 
        \read_value_mux[2][18] , \read_value_mux[2][17] , 
        \read_value_mux[2][16] , \read_value_mux[2][15] , 
        \read_value_mux[2][14] , \read_value_mux[2][13] , 
        \read_value_mux[2][12] , \read_value_mux[2][11] , 
        \read_value_mux[2][10] , \read_value_mux[2][9] , 
        \read_value_mux[2][8] , \read_value_mux[2][7] , \read_value_mux[2][6] , 
        \read_value_mux[2][5] , \read_value_mux[2][4] , \read_value_mux[2][3] , 
        \read_value_mux[2][2] , \read_value_mux[2][1] , \read_value_mux[2][0] , 
        \read_value_mux[1][31] , \read_value_mux[1][30] , 
        \read_value_mux[1][29] , \read_value_mux[1][28] , 
        \read_value_mux[1][27] , \read_value_mux[1][26] , 
        \read_value_mux[1][25] , \read_value_mux[1][24] , 
        \read_value_mux[1][23] , \read_value_mux[1][22] , 
        \read_value_mux[1][21] , \read_value_mux[1][20] , 
        \read_value_mux[1][19] , \read_value_mux[1][18] , 
        \read_value_mux[1][17] , \read_value_mux[1][16] , 
        \read_value_mux[1][15] , \read_value_mux[1][14] , 
        \read_value_mux[1][13] , \read_value_mux[1][12] , 
        \read_value_mux[1][11] , \read_value_mux[1][10] , 
        \read_value_mux[1][9] , \read_value_mux[1][8] , \read_value_mux[1][7] , 
        \read_value_mux[1][6] , \read_value_mux[1][5] , \read_value_mux[1][4] , 
        \read_value_mux[1][3] , \read_value_mux[1][2] , \read_value_mux[1][1] , 
        \read_value_mux[1][0] , \read_value_mux[0][31] , 
        \read_value_mux[0][30] , \read_value_mux[0][29] , 
        \read_value_mux[0][28] , \read_value_mux[0][27] , 
        \read_value_mux[0][26] , \read_value_mux[0][25] , 
        \read_value_mux[0][24] , \read_value_mux[0][23] , 
        \read_value_mux[0][22] , \read_value_mux[0][21] , 
        \read_value_mux[0][20] , \read_value_mux[0][19] , 
        \read_value_mux[0][18] , \read_value_mux[0][17] , 
        \read_value_mux[0][16] , \read_value_mux[0][15] , 
        \read_value_mux[0][14] , \read_value_mux[0][13] , 
        \read_value_mux[0][12] , \read_value_mux[0][11] , 
        \read_value_mux[0][10] , \read_value_mux[0][9] , 
        \read_value_mux[0][8] , \read_value_mux[0][7] , \read_value_mux[0][6] , 
        \read_value_mux[0][5] , \read_value_mux[0][4] , \read_value_mux[0][3] , 
        \read_value_mux[0][2] , \read_value_mux[0][1] , \read_value_mux[0][0] }), .select_i(read_index), .data_o(read_value) );
  DFFX1 \words[31]/data_ff/data_reg[0]  ( .D(\words[31]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[31][0] ) );
  DFFX1 \words[31]/data_ff/data_reg[1]  ( .D(\words[31]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[31][1] ) );
  DFFX1 \words[31]/data_ff/data_reg[2]  ( .D(\words[31]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[31][2] ) );
  DFFX1 \words[31]/data_ff/data_reg[3]  ( .D(\words[31]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[31][3] ), .QN(n1656) );
  DFFX1 \words[31]/data_ff/data_reg[4]  ( .D(\words[31]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[31][4] ) );
  DFFX1 \words[31]/data_ff/data_reg[5]  ( .D(\words[31]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[31][5] ) );
  DFFX1 \words[31]/data_ff/data_reg[6]  ( .D(\words[31]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[31][6] ) );
  DFFX1 \words[31]/data_ff/data_reg[7]  ( .D(\words[31]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[31][7] ) );
  DFFX1 \words[31]/data_ff/data_reg[8]  ( .D(\words[31]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[31][8] ) );
  DFFX1 \words[31]/data_ff/data_reg[9]  ( .D(\words[31]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[31][9] ) );
  DFFX1 \words[31]/data_ff/data_reg[10]  ( .D(\words[31]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[31][10] ) );
  DFFX1 \words[31]/data_ff/data_reg[11]  ( .D(\words[31]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[31][11] ) );
  DFFX1 \words[31]/data_ff/data_reg[12]  ( .D(\words[31]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[31][12] ) );
  DFFX1 \words[31]/data_ff/data_reg[13]  ( .D(\words[31]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[31][13] ) );
  DFFX1 \words[31]/data_ff/data_reg[14]  ( .D(\words[31]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[31][14] ) );
  DFFX1 \words[31]/data_ff/data_reg[15]  ( .D(\words[31]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[31][15] ) );
  DFFX1 \words[31]/data_ff/data_reg[16]  ( .D(\words[31]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[31][16] ) );
  DFFX1 \words[31]/data_ff/data_reg[17]  ( .D(\words[31]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[31][17] ) );
  DFFX1 \words[31]/data_ff/data_reg[18]  ( .D(\words[31]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[31][18] ) );
  DFFX1 \words[31]/data_ff/data_reg[19]  ( .D(\words[31]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[31][19] ) );
  DFFX1 \words[31]/data_ff/data_reg[20]  ( .D(\words[31]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[31][20] ) );
  DFFX1 \words[31]/data_ff/data_reg[21]  ( .D(\words[31]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[31][21] ) );
  DFFX1 \words[31]/data_ff/data_reg[22]  ( .D(\words[31]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[31][22] ) );
  DFFX1 \words[31]/data_ff/data_reg[23]  ( .D(\words[31]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[31][23] ), .QN(n1657) );
  DFFX1 \words[31]/data_ff/data_reg[24]  ( .D(\words[31]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[31][24] ) );
  DFFX1 \words[31]/data_ff/data_reg[25]  ( .D(\words[31]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[31][25] ) );
  DFFX1 \words[31]/data_ff/data_reg[26]  ( .D(\words[31]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[31][26] ) );
  DFFX1 \words[31]/data_ff/data_reg[27]  ( .D(\words[31]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[31][27] ) );
  DFFX1 \words[31]/data_ff/data_reg[28]  ( .D(\words[31]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[31][28] ) );
  DFFX1 \words[31]/data_ff/data_reg[29]  ( .D(\words[31]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[31][29] ) );
  DFFX1 \words[31]/data_ff/data_reg[30]  ( .D(\words[31]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[31][30] ) );
  DFFX1 \words[31]/data_ff/data_reg[31]  ( .D(\words[31]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[31][31] ) );
  DFFX1 \words[31]/valid_ff/data_reg[0]  ( .D(\words[31]/valid_i ), .CLK(clk), 
        .Q(\words[31]/valid_o ) );
  DFFX1 \words[0]/data_ff/data_reg[0]  ( .D(\words[0]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[0][0] ) );
  DFFX1 \words[0]/data_ff/data_reg[1]  ( .D(\words[0]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[0][1] ) );
  DFFX1 \words[0]/data_ff/data_reg[2]  ( .D(\words[0]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[0][2] ) );
  DFFX1 \words[0]/data_ff/data_reg[3]  ( .D(\words[0]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[0][3] ) );
  DFFX1 \words[0]/data_ff/data_reg[4]  ( .D(\words[0]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[0][4] ) );
  DFFX1 \words[0]/data_ff/data_reg[5]  ( .D(\words[0]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[0][5] ) );
  DFFX1 \words[0]/data_ff/data_reg[6]  ( .D(\words[0]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[0][6] ) );
  DFFX1 \words[0]/data_ff/data_reg[7]  ( .D(\words[0]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[0][7] ) );
  DFFX1 \words[0]/data_ff/data_reg[8]  ( .D(\words[0]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[0][8] ) );
  DFFX1 \words[0]/data_ff/data_reg[9]  ( .D(\words[0]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[0][9] ) );
  DFFX1 \words[0]/data_ff/data_reg[10]  ( .D(\words[0]/data_i[10] ), .CLK(clk), 
        .Q(\read_value_mux[0][10] ) );
  DFFX1 \words[0]/data_ff/data_reg[11]  ( .D(\words[0]/data_i[11] ), .CLK(clk), 
        .Q(\read_value_mux[0][11] ) );
  DFFX1 \words[0]/data_ff/data_reg[12]  ( .D(\words[0]/data_i[12] ), .CLK(clk), 
        .Q(\read_value_mux[0][12] ) );
  DFFX1 \words[0]/data_ff/data_reg[13]  ( .D(\words[0]/data_i[13] ), .CLK(clk), 
        .Q(\read_value_mux[0][13] ) );
  DFFX1 \words[0]/data_ff/data_reg[14]  ( .D(\words[0]/data_i[14] ), .CLK(clk), 
        .Q(\read_value_mux[0][14] ) );
  DFFX1 \words[0]/data_ff/data_reg[15]  ( .D(\words[0]/data_i[15] ), .CLK(clk), 
        .Q(\read_value_mux[0][15] ) );
  DFFX1 \words[0]/data_ff/data_reg[16]  ( .D(\words[0]/data_i[16] ), .CLK(clk), 
        .Q(\read_value_mux[0][16] ) );
  DFFX1 \words[0]/data_ff/data_reg[17]  ( .D(\words[0]/data_i[17] ), .CLK(clk), 
        .Q(\read_value_mux[0][17] ) );
  DFFX1 \words[0]/data_ff/data_reg[18]  ( .D(\words[0]/data_i[18] ), .CLK(clk), 
        .Q(\read_value_mux[0][18] ) );
  DFFX1 \words[0]/data_ff/data_reg[19]  ( .D(\words[0]/data_i[19] ), .CLK(clk), 
        .Q(\read_value_mux[0][19] ) );
  DFFX1 \words[0]/data_ff/data_reg[20]  ( .D(\words[0]/data_i[20] ), .CLK(clk), 
        .Q(\read_value_mux[0][20] ) );
  DFFX1 \words[0]/data_ff/data_reg[21]  ( .D(\words[0]/data_i[21] ), .CLK(clk), 
        .Q(\read_value_mux[0][21] ) );
  DFFX1 \words[0]/data_ff/data_reg[22]  ( .D(\words[0]/data_i[22] ), .CLK(clk), 
        .Q(\read_value_mux[0][22] ) );
  DFFX1 \words[0]/data_ff/data_reg[23]  ( .D(\words[0]/data_i[23] ), .CLK(clk), 
        .Q(\read_value_mux[0][23] ) );
  DFFX1 \words[0]/data_ff/data_reg[24]  ( .D(\words[0]/data_i[24] ), .CLK(clk), 
        .Q(\read_value_mux[0][24] ) );
  DFFX1 \words[0]/data_ff/data_reg[25]  ( .D(\words[0]/data_i[25] ), .CLK(clk), 
        .Q(\read_value_mux[0][25] ) );
  DFFX1 \words[0]/data_ff/data_reg[26]  ( .D(\words[0]/data_i[26] ), .CLK(clk), 
        .Q(\read_value_mux[0][26] ) );
  DFFX1 \words[0]/data_ff/data_reg[27]  ( .D(\words[0]/data_i[27] ), .CLK(clk), 
        .Q(\read_value_mux[0][27] ), .QN(n1650) );
  DFFX1 \words[0]/data_ff/data_reg[28]  ( .D(\words[0]/data_i[28] ), .CLK(clk), 
        .Q(\read_value_mux[0][28] ) );
  DFFX1 \words[0]/data_ff/data_reg[29]  ( .D(\words[0]/data_i[29] ), .CLK(clk), 
        .Q(\read_value_mux[0][29] ) );
  DFFX1 \words[0]/data_ff/data_reg[30]  ( .D(\words[0]/data_i[30] ), .CLK(clk), 
        .Q(\read_value_mux[0][30] ) );
  DFFX1 \words[0]/data_ff/data_reg[31]  ( .D(\words[0]/data_i[31] ), .CLK(clk), 
        .Q(\read_value_mux[0][31] ) );
  DFFX1 \words[1]/data_ff/data_reg[0]  ( .D(\words[1]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[1][0] ) );
  DFFX1 \words[1]/data_ff/data_reg[1]  ( .D(\words[1]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[1][1] ) );
  DFFX1 \words[1]/data_ff/data_reg[2]  ( .D(\words[1]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[1][2] ) );
  DFFX1 \words[1]/data_ff/data_reg[3]  ( .D(\words[1]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[1][3] ) );
  DFFX1 \words[1]/data_ff/data_reg[4]  ( .D(\words[1]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[1][4] ) );
  DFFX1 \words[1]/data_ff/data_reg[5]  ( .D(\words[1]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[1][5] ) );
  DFFX1 \words[1]/data_ff/data_reg[6]  ( .D(\words[1]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[1][6] ) );
  DFFX1 \words[1]/data_ff/data_reg[7]  ( .D(\words[1]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[1][7] ) );
  DFFX1 \words[1]/data_ff/data_reg[8]  ( .D(\words[1]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[1][8] ) );
  DFFX1 \words[1]/data_ff/data_reg[9]  ( .D(\words[1]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[1][9] ) );
  DFFX1 \words[1]/data_ff/data_reg[10]  ( .D(\words[1]/data_i[10] ), .CLK(clk), 
        .Q(\read_value_mux[1][10] ) );
  DFFX1 \words[1]/data_ff/data_reg[11]  ( .D(\words[1]/data_i[11] ), .CLK(clk), 
        .Q(\read_value_mux[1][11] ) );
  DFFX1 \words[1]/data_ff/data_reg[12]  ( .D(\words[1]/data_i[12] ), .CLK(clk), 
        .Q(\read_value_mux[1][12] ) );
  DFFX1 \words[1]/data_ff/data_reg[13]  ( .D(\words[1]/data_i[13] ), .CLK(clk), 
        .Q(\read_value_mux[1][13] ) );
  DFFX1 \words[1]/data_ff/data_reg[14]  ( .D(\words[1]/data_i[14] ), .CLK(clk), 
        .Q(\read_value_mux[1][14] ) );
  DFFX1 \words[1]/data_ff/data_reg[15]  ( .D(\words[1]/data_i[15] ), .CLK(clk), 
        .Q(\read_value_mux[1][15] ) );
  DFFX1 \words[1]/data_ff/data_reg[16]  ( .D(\words[1]/data_i[16] ), .CLK(clk), 
        .Q(\read_value_mux[1][16] ) );
  DFFX1 \words[1]/data_ff/data_reg[17]  ( .D(\words[1]/data_i[17] ), .CLK(clk), 
        .Q(\read_value_mux[1][17] ) );
  DFFX1 \words[1]/data_ff/data_reg[18]  ( .D(\words[1]/data_i[18] ), .CLK(clk), 
        .Q(\read_value_mux[1][18] ) );
  DFFX1 \words[1]/data_ff/data_reg[19]  ( .D(\words[1]/data_i[19] ), .CLK(clk), 
        .Q(\read_value_mux[1][19] ) );
  DFFX1 \words[1]/data_ff/data_reg[20]  ( .D(\words[1]/data_i[20] ), .CLK(clk), 
        .Q(\read_value_mux[1][20] ) );
  DFFX1 \words[1]/data_ff/data_reg[21]  ( .D(\words[1]/data_i[21] ), .CLK(clk), 
        .Q(\read_value_mux[1][21] ) );
  DFFX1 \words[1]/data_ff/data_reg[22]  ( .D(\words[1]/data_i[22] ), .CLK(clk), 
        .Q(\read_value_mux[1][22] ) );
  DFFX1 \words[1]/data_ff/data_reg[23]  ( .D(\words[1]/data_i[23] ), .CLK(clk), 
        .Q(\read_value_mux[1][23] ) );
  DFFX1 \words[1]/data_ff/data_reg[24]  ( .D(\words[1]/data_i[24] ), .CLK(clk), 
        .Q(\read_value_mux[1][24] ) );
  DFFX1 \words[1]/data_ff/data_reg[25]  ( .D(\words[1]/data_i[25] ), .CLK(clk), 
        .Q(\read_value_mux[1][25] ) );
  DFFX1 \words[1]/data_ff/data_reg[26]  ( .D(\words[1]/data_i[26] ), .CLK(clk), 
        .Q(\read_value_mux[1][26] ) );
  DFFX1 \words[1]/data_ff/data_reg[27]  ( .D(\words[1]/data_i[27] ), .CLK(clk), 
        .Q(\read_value_mux[1][27] ) );
  DFFX1 \words[1]/data_ff/data_reg[28]  ( .D(\words[1]/data_i[28] ), .CLK(clk), 
        .Q(\read_value_mux[1][28] ) );
  DFFX1 \words[1]/data_ff/data_reg[29]  ( .D(\words[1]/data_i[29] ), .CLK(clk), 
        .Q(\read_value_mux[1][29] ) );
  DFFX1 \words[1]/data_ff/data_reg[30]  ( .D(\words[1]/data_i[30] ), .CLK(clk), 
        .Q(\read_value_mux[1][30] ) );
  DFFX1 \words[1]/data_ff/data_reg[31]  ( .D(\words[1]/data_i[31] ), .CLK(clk), 
        .Q(\read_value_mux[1][31] ) );
  DFFX1 \words[2]/data_ff/data_reg[0]  ( .D(\words[2]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[2][0] ) );
  DFFX1 \words[2]/data_ff/data_reg[1]  ( .D(\words[2]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[2][1] ) );
  DFFX1 \words[2]/data_ff/data_reg[2]  ( .D(\words[2]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[2][2] ) );
  DFFX1 \words[2]/data_ff/data_reg[3]  ( .D(\words[2]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[2][3] ) );
  DFFX1 \words[2]/data_ff/data_reg[4]  ( .D(\words[2]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[2][4] ) );
  DFFX1 \words[2]/data_ff/data_reg[5]  ( .D(\words[2]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[2][5] ), .QN(n1651) );
  DFFX1 \words[2]/data_ff/data_reg[6]  ( .D(\words[2]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[2][6] ) );
  DFFX1 \words[2]/data_ff/data_reg[7]  ( .D(\words[2]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[2][7] ) );
  DFFX1 \words[2]/data_ff/data_reg[8]  ( .D(\words[2]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[2][8] ) );
  DFFX1 \words[2]/data_ff/data_reg[9]  ( .D(\words[2]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[2][9] ) );
  DFFX1 \words[2]/data_ff/data_reg[10]  ( .D(\words[2]/data_i[10] ), .CLK(clk), 
        .Q(\read_value_mux[2][10] ) );
  DFFX1 \words[2]/data_ff/data_reg[11]  ( .D(\words[2]/data_i[11] ), .CLK(clk), 
        .Q(\read_value_mux[2][11] ) );
  DFFX1 \words[2]/data_ff/data_reg[12]  ( .D(\words[2]/data_i[12] ), .CLK(clk), 
        .Q(\read_value_mux[2][12] ) );
  DFFX1 \words[2]/data_ff/data_reg[13]  ( .D(\words[2]/data_i[13] ), .CLK(clk), 
        .Q(\read_value_mux[2][13] ) );
  DFFX1 \words[2]/data_ff/data_reg[14]  ( .D(\words[2]/data_i[14] ), .CLK(clk), 
        .Q(\read_value_mux[2][14] ) );
  DFFX1 \words[2]/data_ff/data_reg[15]  ( .D(\words[2]/data_i[15] ), .CLK(clk), 
        .Q(\read_value_mux[2][15] ) );
  DFFX1 \words[2]/data_ff/data_reg[16]  ( .D(\words[2]/data_i[16] ), .CLK(clk), 
        .Q(\read_value_mux[2][16] ) );
  DFFX1 \words[2]/data_ff/data_reg[17]  ( .D(\words[2]/data_i[17] ), .CLK(clk), 
        .Q(\read_value_mux[2][17] ) );
  DFFX1 \words[2]/data_ff/data_reg[18]  ( .D(\words[2]/data_i[18] ), .CLK(clk), 
        .Q(\read_value_mux[2][18] ) );
  DFFX1 \words[2]/data_ff/data_reg[19]  ( .D(\words[2]/data_i[19] ), .CLK(clk), 
        .Q(\read_value_mux[2][19] ) );
  DFFX1 \words[2]/data_ff/data_reg[20]  ( .D(\words[2]/data_i[20] ), .CLK(clk), 
        .Q(\read_value_mux[2][20] ) );
  DFFX1 \words[2]/data_ff/data_reg[21]  ( .D(\words[2]/data_i[21] ), .CLK(clk), 
        .Q(\read_value_mux[2][21] ) );
  DFFX1 \words[2]/data_ff/data_reg[22]  ( .D(\words[2]/data_i[22] ), .CLK(clk), 
        .Q(\read_value_mux[2][22] ) );
  DFFX1 \words[2]/data_ff/data_reg[23]  ( .D(\words[2]/data_i[23] ), .CLK(clk), 
        .Q(\read_value_mux[2][23] ) );
  DFFX1 \words[2]/data_ff/data_reg[24]  ( .D(\words[2]/data_i[24] ), .CLK(clk), 
        .Q(\read_value_mux[2][24] ) );
  DFFX1 \words[2]/data_ff/data_reg[25]  ( .D(\words[2]/data_i[25] ), .CLK(clk), 
        .Q(\read_value_mux[2][25] ) );
  DFFX1 \words[2]/data_ff/data_reg[26]  ( .D(\words[2]/data_i[26] ), .CLK(clk), 
        .Q(\read_value_mux[2][26] ) );
  DFFX1 \words[2]/data_ff/data_reg[27]  ( .D(\words[2]/data_i[27] ), .CLK(clk), 
        .Q(\read_value_mux[2][27] ) );
  DFFX1 \words[2]/data_ff/data_reg[28]  ( .D(\words[2]/data_i[28] ), .CLK(clk), 
        .Q(\read_value_mux[2][28] ) );
  DFFX1 \words[2]/data_ff/data_reg[29]  ( .D(\words[2]/data_i[29] ), .CLK(clk), 
        .Q(\read_value_mux[2][29] ) );
  DFFX1 \words[2]/data_ff/data_reg[30]  ( .D(\words[2]/data_i[30] ), .CLK(clk), 
        .Q(\read_value_mux[2][30] ) );
  DFFX1 \words[2]/data_ff/data_reg[31]  ( .D(\words[2]/data_i[31] ), .CLK(clk), 
        .Q(\read_value_mux[2][31] ) );
  DFFX1 \words[3]/data_ff/data_reg[0]  ( .D(\words[3]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[3][0] ) );
  DFFX1 \words[3]/data_ff/data_reg[1]  ( .D(\words[3]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[3][1] ) );
  DFFX1 \words[3]/data_ff/data_reg[2]  ( .D(\words[3]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[3][2] ) );
  DFFX1 \words[3]/data_ff/data_reg[3]  ( .D(\words[3]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[3][3] ) );
  DFFX1 \words[3]/data_ff/data_reg[4]  ( .D(\words[3]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[3][4] ) );
  DFFX1 \words[3]/data_ff/data_reg[5]  ( .D(\words[3]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[3][5] ) );
  DFFX1 \words[3]/data_ff/data_reg[6]  ( .D(\words[3]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[3][6] ) );
  DFFX1 \words[3]/data_ff/data_reg[7]  ( .D(\words[3]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[3][7] ) );
  DFFX1 \words[3]/data_ff/data_reg[8]  ( .D(\words[3]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[3][8] ) );
  DFFX1 \words[3]/data_ff/data_reg[9]  ( .D(\words[3]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[3][9] ) );
  DFFX1 \words[3]/data_ff/data_reg[10]  ( .D(\words[3]/data_i[10] ), .CLK(clk), 
        .Q(\read_value_mux[3][10] ) );
  DFFX1 \words[3]/data_ff/data_reg[11]  ( .D(\words[3]/data_i[11] ), .CLK(clk), 
        .Q(\read_value_mux[3][11] ) );
  DFFX1 \words[3]/data_ff/data_reg[12]  ( .D(\words[3]/data_i[12] ), .CLK(clk), 
        .Q(\read_value_mux[3][12] ) );
  DFFX1 \words[3]/data_ff/data_reg[13]  ( .D(\words[3]/data_i[13] ), .CLK(clk), 
        .Q(\read_value_mux[3][13] ) );
  DFFX1 \words[3]/data_ff/data_reg[14]  ( .D(\words[3]/data_i[14] ), .CLK(clk), 
        .Q(\read_value_mux[3][14] ) );
  DFFX1 \words[3]/data_ff/data_reg[15]  ( .D(\words[3]/data_i[15] ), .CLK(clk), 
        .Q(\read_value_mux[3][15] ) );
  DFFX1 \words[3]/data_ff/data_reg[16]  ( .D(\words[3]/data_i[16] ), .CLK(clk), 
        .Q(\read_value_mux[3][16] ) );
  DFFX1 \words[3]/data_ff/data_reg[17]  ( .D(\words[3]/data_i[17] ), .CLK(clk), 
        .Q(\read_value_mux[3][17] ) );
  DFFX1 \words[3]/data_ff/data_reg[18]  ( .D(\words[3]/data_i[18] ), .CLK(clk), 
        .Q(\read_value_mux[3][18] ) );
  DFFX1 \words[3]/data_ff/data_reg[19]  ( .D(\words[3]/data_i[19] ), .CLK(clk), 
        .Q(\read_value_mux[3][19] ) );
  DFFX1 \words[3]/data_ff/data_reg[20]  ( .D(\words[3]/data_i[20] ), .CLK(clk), 
        .Q(\read_value_mux[3][20] ) );
  DFFX1 \words[3]/data_ff/data_reg[21]  ( .D(\words[3]/data_i[21] ), .CLK(clk), 
        .Q(\read_value_mux[3][21] ) );
  DFFX1 \words[3]/data_ff/data_reg[22]  ( .D(\words[3]/data_i[22] ), .CLK(clk), 
        .Q(\read_value_mux[3][22] ) );
  DFFX1 \words[3]/data_ff/data_reg[23]  ( .D(\words[3]/data_i[23] ), .CLK(clk), 
        .Q(\read_value_mux[3][23] ) );
  DFFX1 \words[3]/data_ff/data_reg[24]  ( .D(\words[3]/data_i[24] ), .CLK(clk), 
        .Q(\read_value_mux[3][24] ) );
  DFFX1 \words[3]/data_ff/data_reg[25]  ( .D(\words[3]/data_i[25] ), .CLK(clk), 
        .Q(\read_value_mux[3][25] ) );
  DFFX1 \words[3]/data_ff/data_reg[26]  ( .D(\words[3]/data_i[26] ), .CLK(clk), 
        .Q(\read_value_mux[3][26] ) );
  DFFX1 \words[3]/data_ff/data_reg[27]  ( .D(\words[3]/data_i[27] ), .CLK(clk), 
        .Q(\read_value_mux[3][27] ) );
  DFFX1 \words[3]/data_ff/data_reg[28]  ( .D(\words[3]/data_i[28] ), .CLK(clk), 
        .Q(\read_value_mux[3][28] ) );
  DFFX1 \words[3]/data_ff/data_reg[29]  ( .D(\words[3]/data_i[29] ), .CLK(clk), 
        .Q(\read_value_mux[3][29] ) );
  DFFX1 \words[3]/data_ff/data_reg[30]  ( .D(\words[3]/data_i[30] ), .CLK(clk), 
        .Q(\read_value_mux[3][30] ) );
  DFFX1 \words[3]/data_ff/data_reg[31]  ( .D(\words[3]/data_i[31] ), .CLK(clk), 
        .Q(\read_value_mux[3][31] ) );
  DFFX1 \words[4]/data_ff/data_reg[0]  ( .D(\words[4]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[4][0] ) );
  DFFX1 \words[4]/data_ff/data_reg[1]  ( .D(\words[4]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[4][1] ) );
  DFFX1 \words[4]/data_ff/data_reg[2]  ( .D(\words[4]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[4][2] ) );
  DFFX1 \words[4]/data_ff/data_reg[3]  ( .D(\words[4]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[4][3] ) );
  DFFX1 \words[4]/data_ff/data_reg[4]  ( .D(\words[4]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[4][4] ) );
  DFFX1 \words[4]/data_ff/data_reg[5]  ( .D(\words[4]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[4][5] ) );
  DFFX1 \words[4]/data_ff/data_reg[6]  ( .D(\words[4]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[4][6] ) );
  DFFX1 \words[4]/data_ff/data_reg[7]  ( .D(\words[4]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[4][7] ) );
  DFFX1 \words[4]/data_ff/data_reg[8]  ( .D(\words[4]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[4][8] ) );
  DFFX1 \words[4]/data_ff/data_reg[9]  ( .D(\words[4]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[4][9] ) );
  DFFX1 \words[4]/data_ff/data_reg[10]  ( .D(\words[4]/data_i[10] ), .CLK(clk), 
        .Q(\read_value_mux[4][10] ) );
  DFFX1 \words[4]/data_ff/data_reg[11]  ( .D(\words[4]/data_i[11] ), .CLK(clk), 
        .Q(\read_value_mux[4][11] ) );
  DFFX1 \words[4]/data_ff/data_reg[12]  ( .D(\words[4]/data_i[12] ), .CLK(clk), 
        .Q(\read_value_mux[4][12] ) );
  DFFX1 \words[4]/data_ff/data_reg[13]  ( .D(\words[4]/data_i[13] ), .CLK(clk), 
        .Q(\read_value_mux[4][13] ) );
  DFFX1 \words[4]/data_ff/data_reg[14]  ( .D(\words[4]/data_i[14] ), .CLK(clk), 
        .Q(\read_value_mux[4][14] ) );
  DFFX1 \words[4]/data_ff/data_reg[15]  ( .D(\words[4]/data_i[15] ), .CLK(clk), 
        .Q(\read_value_mux[4][15] ) );
  DFFX1 \words[4]/data_ff/data_reg[16]  ( .D(\words[4]/data_i[16] ), .CLK(clk), 
        .Q(\read_value_mux[4][16] ) );
  DFFX1 \words[4]/data_ff/data_reg[17]  ( .D(\words[4]/data_i[17] ), .CLK(clk), 
        .Q(\read_value_mux[4][17] ) );
  DFFX1 \words[4]/data_ff/data_reg[18]  ( .D(\words[4]/data_i[18] ), .CLK(clk), 
        .Q(\read_value_mux[4][18] ) );
  DFFX1 \words[4]/data_ff/data_reg[19]  ( .D(\words[4]/data_i[19] ), .CLK(clk), 
        .Q(\read_value_mux[4][19] ) );
  DFFX1 \words[4]/data_ff/data_reg[20]  ( .D(\words[4]/data_i[20] ), .CLK(clk), 
        .Q(\read_value_mux[4][20] ) );
  DFFX1 \words[4]/data_ff/data_reg[21]  ( .D(\words[4]/data_i[21] ), .CLK(clk), 
        .Q(\read_value_mux[4][21] ) );
  DFFX1 \words[4]/data_ff/data_reg[22]  ( .D(\words[4]/data_i[22] ), .CLK(clk), 
        .Q(\read_value_mux[4][22] ) );
  DFFX1 \words[4]/data_ff/data_reg[23]  ( .D(\words[4]/data_i[23] ), .CLK(clk), 
        .Q(\read_value_mux[4][23] ) );
  DFFX1 \words[4]/data_ff/data_reg[24]  ( .D(\words[4]/data_i[24] ), .CLK(clk), 
        .Q(\read_value_mux[4][24] ) );
  DFFX1 \words[4]/data_ff/data_reg[25]  ( .D(\words[4]/data_i[25] ), .CLK(clk), 
        .Q(\read_value_mux[4][25] ) );
  DFFX1 \words[4]/data_ff/data_reg[26]  ( .D(\words[4]/data_i[26] ), .CLK(clk), 
        .Q(\read_value_mux[4][26] ) );
  DFFX1 \words[4]/data_ff/data_reg[27]  ( .D(\words[4]/data_i[27] ), .CLK(clk), 
        .Q(\read_value_mux[4][27] ) );
  DFFX1 \words[4]/data_ff/data_reg[28]  ( .D(\words[4]/data_i[28] ), .CLK(clk), 
        .Q(\read_value_mux[4][28] ) );
  DFFX1 \words[4]/data_ff/data_reg[29]  ( .D(\words[4]/data_i[29] ), .CLK(clk), 
        .Q(\read_value_mux[4][29] ) );
  DFFX1 \words[4]/data_ff/data_reg[30]  ( .D(\words[4]/data_i[30] ), .CLK(clk), 
        .Q(\read_value_mux[4][30] ) );
  DFFX1 \words[4]/data_ff/data_reg[31]  ( .D(\words[4]/data_i[31] ), .CLK(clk), 
        .Q(\read_value_mux[4][31] ) );
  DFFX1 \words[5]/data_ff/data_reg[0]  ( .D(\words[5]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[5][0] ) );
  DFFX1 \words[5]/data_ff/data_reg[1]  ( .D(\words[5]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[5][1] ) );
  DFFX1 \words[5]/data_ff/data_reg[2]  ( .D(\words[5]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[5][2] ) );
  DFFX1 \words[5]/data_ff/data_reg[3]  ( .D(\words[5]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[5][3] ) );
  DFFX1 \words[5]/data_ff/data_reg[4]  ( .D(\words[5]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[5][4] ) );
  DFFX1 \words[5]/data_ff/data_reg[5]  ( .D(\words[5]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[5][5] ) );
  DFFX1 \words[5]/data_ff/data_reg[6]  ( .D(\words[5]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[5][6] ) );
  DFFX1 \words[5]/data_ff/data_reg[7]  ( .D(\words[5]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[5][7] ) );
  DFFX1 \words[5]/data_ff/data_reg[8]  ( .D(\words[5]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[5][8] ) );
  DFFX1 \words[5]/data_ff/data_reg[9]  ( .D(\words[5]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[5][9] ) );
  DFFX1 \words[5]/data_ff/data_reg[10]  ( .D(\words[5]/data_i[10] ), .CLK(clk), 
        .Q(\read_value_mux[5][10] ) );
  DFFX1 \words[5]/data_ff/data_reg[11]  ( .D(\words[5]/data_i[11] ), .CLK(clk), 
        .Q(\read_value_mux[5][11] ) );
  DFFX1 \words[5]/data_ff/data_reg[12]  ( .D(\words[5]/data_i[12] ), .CLK(clk), 
        .Q(\read_value_mux[5][12] ) );
  DFFX1 \words[5]/data_ff/data_reg[13]  ( .D(\words[5]/data_i[13] ), .CLK(clk), 
        .Q(\read_value_mux[5][13] ) );
  DFFX1 \words[5]/data_ff/data_reg[14]  ( .D(\words[5]/data_i[14] ), .CLK(clk), 
        .Q(\read_value_mux[5][14] ) );
  DFFX1 \words[5]/data_ff/data_reg[15]  ( .D(\words[5]/data_i[15] ), .CLK(clk), 
        .Q(\read_value_mux[5][15] ) );
  DFFX1 \words[5]/data_ff/data_reg[16]  ( .D(\words[5]/data_i[16] ), .CLK(clk), 
        .Q(\read_value_mux[5][16] ) );
  DFFX1 \words[5]/data_ff/data_reg[17]  ( .D(\words[5]/data_i[17] ), .CLK(clk), 
        .Q(\read_value_mux[5][17] ) );
  DFFX1 \words[5]/data_ff/data_reg[18]  ( .D(\words[5]/data_i[18] ), .CLK(clk), 
        .Q(\read_value_mux[5][18] ) );
  DFFX1 \words[5]/data_ff/data_reg[19]  ( .D(\words[5]/data_i[19] ), .CLK(clk), 
        .Q(\read_value_mux[5][19] ) );
  DFFX1 \words[5]/data_ff/data_reg[20]  ( .D(\words[5]/data_i[20] ), .CLK(clk), 
        .Q(\read_value_mux[5][20] ) );
  DFFX1 \words[5]/data_ff/data_reg[21]  ( .D(\words[5]/data_i[21] ), .CLK(clk), 
        .Q(\read_value_mux[5][21] ) );
  DFFX1 \words[5]/data_ff/data_reg[22]  ( .D(\words[5]/data_i[22] ), .CLK(clk), 
        .Q(\read_value_mux[5][22] ) );
  DFFX1 \words[5]/data_ff/data_reg[23]  ( .D(\words[5]/data_i[23] ), .CLK(clk), 
        .Q(\read_value_mux[5][23] ) );
  DFFX1 \words[5]/data_ff/data_reg[24]  ( .D(\words[5]/data_i[24] ), .CLK(clk), 
        .Q(\read_value_mux[5][24] ) );
  DFFX1 \words[5]/data_ff/data_reg[25]  ( .D(\words[5]/data_i[25] ), .CLK(clk), 
        .Q(\read_value_mux[5][25] ) );
  DFFX1 \words[5]/data_ff/data_reg[26]  ( .D(\words[5]/data_i[26] ), .CLK(clk), 
        .Q(\read_value_mux[5][26] ) );
  DFFX1 \words[5]/data_ff/data_reg[27]  ( .D(\words[5]/data_i[27] ), .CLK(clk), 
        .Q(\read_value_mux[5][27] ) );
  DFFX1 \words[5]/data_ff/data_reg[28]  ( .D(\words[5]/data_i[28] ), .CLK(clk), 
        .Q(\read_value_mux[5][28] ) );
  DFFX1 \words[5]/data_ff/data_reg[29]  ( .D(\words[5]/data_i[29] ), .CLK(clk), 
        .Q(\read_value_mux[5][29] ) );
  DFFX1 \words[5]/data_ff/data_reg[30]  ( .D(\words[5]/data_i[30] ), .CLK(clk), 
        .Q(\read_value_mux[5][30] ) );
  DFFX1 \words[5]/data_ff/data_reg[31]  ( .D(\words[5]/data_i[31] ), .CLK(clk), 
        .Q(\read_value_mux[5][31] ) );
  DFFX1 \words[6]/data_ff/data_reg[0]  ( .D(\words[6]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[6][0] ) );
  DFFX1 \words[6]/data_ff/data_reg[1]  ( .D(\words[6]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[6][1] ) );
  DFFX1 \words[6]/data_ff/data_reg[2]  ( .D(\words[6]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[6][2] ) );
  DFFX1 \words[6]/data_ff/data_reg[3]  ( .D(\words[6]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[6][3] ) );
  DFFX1 \words[6]/data_ff/data_reg[4]  ( .D(\words[6]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[6][4] ) );
  DFFX1 \words[6]/data_ff/data_reg[5]  ( .D(\words[6]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[6][5] ) );
  DFFX1 \words[6]/data_ff/data_reg[6]  ( .D(\words[6]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[6][6] ) );
  DFFX1 \words[6]/data_ff/data_reg[7]  ( .D(\words[6]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[6][7] ) );
  DFFX1 \words[6]/data_ff/data_reg[8]  ( .D(\words[6]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[6][8] ) );
  DFFX1 \words[6]/data_ff/data_reg[9]  ( .D(\words[6]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[6][9] ) );
  DFFX1 \words[6]/data_ff/data_reg[10]  ( .D(\words[6]/data_i[10] ), .CLK(clk), 
        .Q(\read_value_mux[6][10] ) );
  DFFX1 \words[6]/data_ff/data_reg[11]  ( .D(\words[6]/data_i[11] ), .CLK(clk), 
        .Q(\read_value_mux[6][11] ) );
  DFFX1 \words[6]/data_ff/data_reg[12]  ( .D(\words[6]/data_i[12] ), .CLK(clk), 
        .Q(\read_value_mux[6][12] ) );
  DFFX1 \words[6]/data_ff/data_reg[13]  ( .D(\words[6]/data_i[13] ), .CLK(clk), 
        .Q(\read_value_mux[6][13] ) );
  DFFX1 \words[6]/data_ff/data_reg[14]  ( .D(\words[6]/data_i[14] ), .CLK(clk), 
        .Q(\read_value_mux[6][14] ) );
  DFFX1 \words[6]/data_ff/data_reg[15]  ( .D(\words[6]/data_i[15] ), .CLK(clk), 
        .Q(\read_value_mux[6][15] ) );
  DFFX1 \words[6]/data_ff/data_reg[16]  ( .D(\words[6]/data_i[16] ), .CLK(clk), 
        .Q(\read_value_mux[6][16] ) );
  DFFX1 \words[6]/data_ff/data_reg[17]  ( .D(\words[6]/data_i[17] ), .CLK(clk), 
        .Q(\read_value_mux[6][17] ) );
  DFFX1 \words[6]/data_ff/data_reg[18]  ( .D(\words[6]/data_i[18] ), .CLK(clk), 
        .Q(\read_value_mux[6][18] ) );
  DFFX1 \words[6]/data_ff/data_reg[19]  ( .D(\words[6]/data_i[19] ), .CLK(clk), 
        .Q(\read_value_mux[6][19] ) );
  DFFX1 \words[6]/data_ff/data_reg[20]  ( .D(\words[6]/data_i[20] ), .CLK(clk), 
        .Q(\read_value_mux[6][20] ) );
  DFFX1 \words[6]/data_ff/data_reg[21]  ( .D(\words[6]/data_i[21] ), .CLK(clk), 
        .Q(\read_value_mux[6][21] ) );
  DFFX1 \words[6]/data_ff/data_reg[22]  ( .D(\words[6]/data_i[22] ), .CLK(clk), 
        .Q(\read_value_mux[6][22] ) );
  DFFX1 \words[6]/data_ff/data_reg[23]  ( .D(\words[6]/data_i[23] ), .CLK(clk), 
        .Q(\read_value_mux[6][23] ) );
  DFFX1 \words[6]/data_ff/data_reg[24]  ( .D(\words[6]/data_i[24] ), .CLK(clk), 
        .Q(\read_value_mux[6][24] ) );
  DFFX1 \words[6]/data_ff/data_reg[25]  ( .D(\words[6]/data_i[25] ), .CLK(clk), 
        .Q(\read_value_mux[6][25] ) );
  DFFX1 \words[6]/data_ff/data_reg[26]  ( .D(\words[6]/data_i[26] ), .CLK(clk), 
        .Q(\read_value_mux[6][26] ) );
  DFFX1 \words[6]/data_ff/data_reg[27]  ( .D(\words[6]/data_i[27] ), .CLK(clk), 
        .Q(\read_value_mux[6][27] ) );
  DFFX1 \words[6]/data_ff/data_reg[28]  ( .D(\words[6]/data_i[28] ), .CLK(clk), 
        .Q(\read_value_mux[6][28] ) );
  DFFX1 \words[6]/data_ff/data_reg[29]  ( .D(\words[6]/data_i[29] ), .CLK(clk), 
        .Q(\read_value_mux[6][29] ) );
  DFFX1 \words[6]/data_ff/data_reg[30]  ( .D(\words[6]/data_i[30] ), .CLK(clk), 
        .Q(\read_value_mux[6][30] ) );
  DFFX1 \words[6]/data_ff/data_reg[31]  ( .D(\words[6]/data_i[31] ), .CLK(clk), 
        .Q(\read_value_mux[6][31] ) );
  DFFX1 \words[7]/data_ff/data_reg[0]  ( .D(\words[7]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[7][0] ) );
  DFFX1 \words[7]/data_ff/data_reg[1]  ( .D(\words[7]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[7][1] ) );
  DFFX1 \words[7]/data_ff/data_reg[2]  ( .D(\words[7]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[7][2] ) );
  DFFX1 \words[7]/data_ff/data_reg[3]  ( .D(\words[7]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[7][3] ) );
  DFFX1 \words[7]/data_ff/data_reg[4]  ( .D(\words[7]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[7][4] ) );
  DFFX1 \words[7]/data_ff/data_reg[5]  ( .D(\words[7]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[7][5] ) );
  DFFX1 \words[7]/data_ff/data_reg[6]  ( .D(\words[7]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[7][6] ) );
  DFFX1 \words[7]/data_ff/data_reg[7]  ( .D(\words[7]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[7][7] ) );
  DFFX1 \words[7]/data_ff/data_reg[8]  ( .D(\words[7]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[7][8] ) );
  DFFX1 \words[7]/data_ff/data_reg[9]  ( .D(\words[7]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[7][9] ) );
  DFFX1 \words[7]/data_ff/data_reg[10]  ( .D(\words[7]/data_i[10] ), .CLK(clk), 
        .Q(\read_value_mux[7][10] ) );
  DFFX1 \words[7]/data_ff/data_reg[11]  ( .D(\words[7]/data_i[11] ), .CLK(clk), 
        .Q(\read_value_mux[7][11] ) );
  DFFX1 \words[7]/data_ff/data_reg[12]  ( .D(\words[7]/data_i[12] ), .CLK(clk), 
        .Q(\read_value_mux[7][12] ) );
  DFFX1 \words[7]/data_ff/data_reg[13]  ( .D(\words[7]/data_i[13] ), .CLK(clk), 
        .Q(\read_value_mux[7][13] ) );
  DFFX1 \words[7]/data_ff/data_reg[14]  ( .D(\words[7]/data_i[14] ), .CLK(clk), 
        .Q(\read_value_mux[7][14] ) );
  DFFX1 \words[7]/data_ff/data_reg[15]  ( .D(\words[7]/data_i[15] ), .CLK(clk), 
        .Q(\read_value_mux[7][15] ) );
  DFFX1 \words[7]/data_ff/data_reg[16]  ( .D(\words[7]/data_i[16] ), .CLK(clk), 
        .Q(\read_value_mux[7][16] ) );
  DFFX1 \words[7]/data_ff/data_reg[17]  ( .D(\words[7]/data_i[17] ), .CLK(clk), 
        .Q(\read_value_mux[7][17] ) );
  DFFX1 \words[7]/data_ff/data_reg[18]  ( .D(\words[7]/data_i[18] ), .CLK(clk), 
        .Q(\read_value_mux[7][18] ) );
  DFFX1 \words[7]/data_ff/data_reg[19]  ( .D(\words[7]/data_i[19] ), .CLK(clk), 
        .Q(\read_value_mux[7][19] ) );
  DFFX1 \words[7]/data_ff/data_reg[20]  ( .D(\words[7]/data_i[20] ), .CLK(clk), 
        .Q(\read_value_mux[7][20] ) );
  DFFX1 \words[7]/data_ff/data_reg[21]  ( .D(\words[7]/data_i[21] ), .CLK(clk), 
        .Q(\read_value_mux[7][21] ) );
  DFFX1 \words[7]/data_ff/data_reg[22]  ( .D(\words[7]/data_i[22] ), .CLK(clk), 
        .Q(\read_value_mux[7][22] ) );
  DFFX1 \words[7]/data_ff/data_reg[23]  ( .D(\words[7]/data_i[23] ), .CLK(clk), 
        .Q(\read_value_mux[7][23] ) );
  DFFX1 \words[7]/data_ff/data_reg[24]  ( .D(\words[7]/data_i[24] ), .CLK(clk), 
        .Q(\read_value_mux[7][24] ) );
  DFFX1 \words[7]/data_ff/data_reg[25]  ( .D(\words[7]/data_i[25] ), .CLK(clk), 
        .Q(\read_value_mux[7][25] ) );
  DFFX1 \words[7]/data_ff/data_reg[26]  ( .D(\words[7]/data_i[26] ), .CLK(clk), 
        .Q(\read_value_mux[7][26] ) );
  DFFX1 \words[7]/data_ff/data_reg[27]  ( .D(\words[7]/data_i[27] ), .CLK(clk), 
        .Q(\read_value_mux[7][27] ) );
  DFFX1 \words[7]/data_ff/data_reg[28]  ( .D(\words[7]/data_i[28] ), .CLK(clk), 
        .Q(\read_value_mux[7][28] ) );
  DFFX1 \words[7]/data_ff/data_reg[29]  ( .D(\words[7]/data_i[29] ), .CLK(clk), 
        .Q(\read_value_mux[7][29] ) );
  DFFX1 \words[7]/data_ff/data_reg[30]  ( .D(\words[7]/data_i[30] ), .CLK(clk), 
        .Q(\read_value_mux[7][30] ) );
  DFFX1 \words[7]/data_ff/data_reg[31]  ( .D(\words[7]/data_i[31] ), .CLK(clk), 
        .Q(\read_value_mux[7][31] ) );
  DFFX1 \words[8]/data_ff/data_reg[0]  ( .D(\words[8]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[8][0] ) );
  DFFX1 \words[8]/data_ff/data_reg[1]  ( .D(\words[8]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[8][1] ) );
  DFFX1 \words[8]/data_ff/data_reg[2]  ( .D(\words[8]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[8][2] ) );
  DFFX1 \words[8]/data_ff/data_reg[3]  ( .D(\words[8]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[8][3] ) );
  DFFX1 \words[8]/data_ff/data_reg[4]  ( .D(\words[8]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[8][4] ) );
  DFFX1 \words[8]/data_ff/data_reg[5]  ( .D(\words[8]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[8][5] ) );
  DFFX1 \words[8]/data_ff/data_reg[6]  ( .D(\words[8]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[8][6] ) );
  DFFX1 \words[8]/data_ff/data_reg[7]  ( .D(\words[8]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[8][7] ) );
  DFFX1 \words[8]/data_ff/data_reg[8]  ( .D(\words[8]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[8][8] ) );
  DFFX1 \words[8]/data_ff/data_reg[9]  ( .D(\words[8]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[8][9] ) );
  DFFX1 \words[8]/data_ff/data_reg[10]  ( .D(\words[8]/data_i[10] ), .CLK(clk), 
        .Q(\read_value_mux[8][10] ) );
  DFFX1 \words[8]/data_ff/data_reg[11]  ( .D(\words[8]/data_i[11] ), .CLK(clk), 
        .Q(\read_value_mux[8][11] ) );
  DFFX1 \words[8]/data_ff/data_reg[12]  ( .D(\words[8]/data_i[12] ), .CLK(clk), 
        .Q(\read_value_mux[8][12] ) );
  DFFX1 \words[8]/data_ff/data_reg[13]  ( .D(\words[8]/data_i[13] ), .CLK(clk), 
        .Q(\read_value_mux[8][13] ) );
  DFFX1 \words[8]/data_ff/data_reg[14]  ( .D(\words[8]/data_i[14] ), .CLK(clk), 
        .Q(\read_value_mux[8][14] ) );
  DFFX1 \words[8]/data_ff/data_reg[15]  ( .D(\words[8]/data_i[15] ), .CLK(clk), 
        .Q(\read_value_mux[8][15] ) );
  DFFX1 \words[8]/data_ff/data_reg[16]  ( .D(\words[8]/data_i[16] ), .CLK(clk), 
        .Q(\read_value_mux[8][16] ) );
  DFFX1 \words[8]/data_ff/data_reg[17]  ( .D(\words[8]/data_i[17] ), .CLK(clk), 
        .Q(\read_value_mux[8][17] ) );
  DFFX1 \words[8]/data_ff/data_reg[18]  ( .D(\words[8]/data_i[18] ), .CLK(clk), 
        .Q(\read_value_mux[8][18] ) );
  DFFX1 \words[8]/data_ff/data_reg[19]  ( .D(\words[8]/data_i[19] ), .CLK(clk), 
        .Q(\read_value_mux[8][19] ) );
  DFFX1 \words[8]/data_ff/data_reg[20]  ( .D(\words[8]/data_i[20] ), .CLK(clk), 
        .Q(\read_value_mux[8][20] ) );
  DFFX1 \words[8]/data_ff/data_reg[21]  ( .D(\words[8]/data_i[21] ), .CLK(clk), 
        .Q(\read_value_mux[8][21] ) );
  DFFX1 \words[8]/data_ff/data_reg[22]  ( .D(\words[8]/data_i[22] ), .CLK(clk), 
        .Q(\read_value_mux[8][22] ) );
  DFFX1 \words[8]/data_ff/data_reg[23]  ( .D(\words[8]/data_i[23] ), .CLK(clk), 
        .Q(\read_value_mux[8][23] ) );
  DFFX1 \words[8]/data_ff/data_reg[24]  ( .D(\words[8]/data_i[24] ), .CLK(clk), 
        .Q(\read_value_mux[8][24] ) );
  DFFX1 \words[8]/data_ff/data_reg[25]  ( .D(\words[8]/data_i[25] ), .CLK(clk), 
        .Q(\read_value_mux[8][25] ) );
  DFFX1 \words[8]/data_ff/data_reg[26]  ( .D(\words[8]/data_i[26] ), .CLK(clk), 
        .Q(\read_value_mux[8][26] ) );
  DFFX1 \words[8]/data_ff/data_reg[27]  ( .D(\words[8]/data_i[27] ), .CLK(clk), 
        .Q(\read_value_mux[8][27] ) );
  DFFX1 \words[8]/data_ff/data_reg[28]  ( .D(\words[8]/data_i[28] ), .CLK(clk), 
        .Q(\read_value_mux[8][28] ) );
  DFFX1 \words[8]/data_ff/data_reg[29]  ( .D(\words[8]/data_i[29] ), .CLK(clk), 
        .Q(\read_value_mux[8][29] ) );
  DFFX1 \words[8]/data_ff/data_reg[30]  ( .D(\words[8]/data_i[30] ), .CLK(clk), 
        .Q(\read_value_mux[8][30] ) );
  DFFX1 \words[8]/data_ff/data_reg[31]  ( .D(\words[8]/data_i[31] ), .CLK(clk), 
        .Q(\read_value_mux[8][31] ) );
  DFFX1 \words[9]/data_ff/data_reg[0]  ( .D(\words[9]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[9][0] ) );
  DFFX1 \words[9]/data_ff/data_reg[1]  ( .D(\words[9]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[9][1] ) );
  DFFX1 \words[9]/data_ff/data_reg[2]  ( .D(\words[9]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[9][2] ) );
  DFFX1 \words[9]/data_ff/data_reg[3]  ( .D(\words[9]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[9][3] ) );
  DFFX1 \words[9]/data_ff/data_reg[4]  ( .D(\words[9]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[9][4] ) );
  DFFX1 \words[9]/data_ff/data_reg[5]  ( .D(\words[9]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[9][5] ) );
  DFFX1 \words[9]/data_ff/data_reg[6]  ( .D(\words[9]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[9][6] ) );
  DFFX1 \words[9]/data_ff/data_reg[7]  ( .D(\words[9]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[9][7] ) );
  DFFX1 \words[9]/data_ff/data_reg[8]  ( .D(\words[9]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[9][8] ) );
  DFFX1 \words[9]/data_ff/data_reg[9]  ( .D(\words[9]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[9][9] ) );
  DFFX1 \words[9]/data_ff/data_reg[10]  ( .D(\words[9]/data_i[10] ), .CLK(clk), 
        .Q(\read_value_mux[9][10] ) );
  DFFX1 \words[9]/data_ff/data_reg[11]  ( .D(\words[9]/data_i[11] ), .CLK(clk), 
        .Q(\read_value_mux[9][11] ) );
  DFFX1 \words[9]/data_ff/data_reg[12]  ( .D(\words[9]/data_i[12] ), .CLK(clk), 
        .Q(\read_value_mux[9][12] ) );
  DFFX1 \words[9]/data_ff/data_reg[13]  ( .D(\words[9]/data_i[13] ), .CLK(clk), 
        .Q(\read_value_mux[9][13] ) );
  DFFX1 \words[9]/data_ff/data_reg[14]  ( .D(\words[9]/data_i[14] ), .CLK(clk), 
        .Q(\read_value_mux[9][14] ) );
  DFFX1 \words[9]/data_ff/data_reg[15]  ( .D(\words[9]/data_i[15] ), .CLK(clk), 
        .Q(\read_value_mux[9][15] ) );
  DFFX1 \words[9]/data_ff/data_reg[16]  ( .D(\words[9]/data_i[16] ), .CLK(clk), 
        .Q(\read_value_mux[9][16] ) );
  DFFX1 \words[9]/data_ff/data_reg[17]  ( .D(\words[9]/data_i[17] ), .CLK(clk), 
        .Q(\read_value_mux[9][17] ) );
  DFFX1 \words[9]/data_ff/data_reg[18]  ( .D(\words[9]/data_i[18] ), .CLK(clk), 
        .Q(\read_value_mux[9][18] ) );
  DFFX1 \words[9]/data_ff/data_reg[19]  ( .D(\words[9]/data_i[19] ), .CLK(clk), 
        .Q(\read_value_mux[9][19] ) );
  DFFX1 \words[9]/data_ff/data_reg[20]  ( .D(\words[9]/data_i[20] ), .CLK(clk), 
        .Q(\read_value_mux[9][20] ) );
  DFFX1 \words[9]/data_ff/data_reg[21]  ( .D(\words[9]/data_i[21] ), .CLK(clk), 
        .Q(\read_value_mux[9][21] ) );
  DFFX1 \words[9]/data_ff/data_reg[22]  ( .D(\words[9]/data_i[22] ), .CLK(clk), 
        .Q(\read_value_mux[9][22] ) );
  DFFX1 \words[9]/data_ff/data_reg[23]  ( .D(\words[9]/data_i[23] ), .CLK(clk), 
        .Q(\read_value_mux[9][23] ) );
  DFFX1 \words[9]/data_ff/data_reg[24]  ( .D(\words[9]/data_i[24] ), .CLK(clk), 
        .Q(\read_value_mux[9][24] ) );
  DFFX1 \words[9]/data_ff/data_reg[25]  ( .D(\words[9]/data_i[25] ), .CLK(clk), 
        .Q(\read_value_mux[9][25] ) );
  DFFX1 \words[9]/data_ff/data_reg[26]  ( .D(\words[9]/data_i[26] ), .CLK(clk), 
        .Q(\read_value_mux[9][26] ) );
  DFFX1 \words[9]/data_ff/data_reg[27]  ( .D(\words[9]/data_i[27] ), .CLK(clk), 
        .Q(\read_value_mux[9][27] ) );
  DFFX1 \words[9]/data_ff/data_reg[28]  ( .D(\words[9]/data_i[28] ), .CLK(clk), 
        .Q(\read_value_mux[9][28] ) );
  DFFX1 \words[9]/data_ff/data_reg[29]  ( .D(\words[9]/data_i[29] ), .CLK(clk), 
        .Q(\read_value_mux[9][29] ) );
  DFFX1 \words[9]/data_ff/data_reg[30]  ( .D(\words[9]/data_i[30] ), .CLK(clk), 
        .Q(\read_value_mux[9][30] ) );
  DFFX1 \words[9]/data_ff/data_reg[31]  ( .D(\words[9]/data_i[31] ), .CLK(clk), 
        .Q(\read_value_mux[9][31] ) );
  DFFX1 \words[10]/data_ff/data_reg[0]  ( .D(\words[10]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[10][0] ) );
  DFFX1 \words[10]/data_ff/data_reg[1]  ( .D(\words[10]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[10][1] ) );
  DFFX1 \words[10]/data_ff/data_reg[2]  ( .D(\words[10]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[10][2] ) );
  DFFX1 \words[10]/data_ff/data_reg[3]  ( .D(\words[10]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[10][3] ) );
  DFFX1 \words[10]/data_ff/data_reg[4]  ( .D(\words[10]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[10][4] ) );
  DFFX1 \words[10]/data_ff/data_reg[5]  ( .D(\words[10]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[10][5] ) );
  DFFX1 \words[10]/data_ff/data_reg[6]  ( .D(\words[10]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[10][6] ) );
  DFFX1 \words[10]/data_ff/data_reg[7]  ( .D(\words[10]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[10][7] ) );
  DFFX1 \words[10]/data_ff/data_reg[8]  ( .D(\words[10]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[10][8] ) );
  DFFX1 \words[10]/data_ff/data_reg[9]  ( .D(\words[10]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[10][9] ) );
  DFFX1 \words[10]/data_ff/data_reg[10]  ( .D(\words[10]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[10][10] ) );
  DFFX1 \words[10]/data_ff/data_reg[11]  ( .D(\words[10]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[10][11] ) );
  DFFX1 \words[10]/data_ff/data_reg[12]  ( .D(\words[10]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[10][12] ) );
  DFFX1 \words[10]/data_ff/data_reg[13]  ( .D(\words[10]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[10][13] ) );
  DFFX1 \words[10]/data_ff/data_reg[14]  ( .D(\words[10]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[10][14] ) );
  DFFX1 \words[10]/data_ff/data_reg[15]  ( .D(\words[10]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[10][15] ) );
  DFFX1 \words[10]/data_ff/data_reg[16]  ( .D(\words[10]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[10][16] ) );
  DFFX1 \words[10]/data_ff/data_reg[17]  ( .D(\words[10]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[10][17] ) );
  DFFX1 \words[10]/data_ff/data_reg[18]  ( .D(\words[10]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[10][18] ) );
  DFFX1 \words[10]/data_ff/data_reg[19]  ( .D(\words[10]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[10][19] ) );
  DFFX1 \words[10]/data_ff/data_reg[20]  ( .D(\words[10]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[10][20] ) );
  DFFX1 \words[10]/data_ff/data_reg[21]  ( .D(\words[10]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[10][21] ) );
  DFFX1 \words[10]/data_ff/data_reg[22]  ( .D(\words[10]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[10][22] ) );
  DFFX1 \words[10]/data_ff/data_reg[23]  ( .D(\words[10]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[10][23] ) );
  DFFX1 \words[10]/data_ff/data_reg[24]  ( .D(\words[10]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[10][24] ) );
  DFFX1 \words[10]/data_ff/data_reg[25]  ( .D(\words[10]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[10][25] ) );
  DFFX1 \words[10]/data_ff/data_reg[26]  ( .D(\words[10]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[10][26] ) );
  DFFX1 \words[10]/data_ff/data_reg[27]  ( .D(\words[10]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[10][27] ) );
  DFFX1 \words[10]/data_ff/data_reg[28]  ( .D(\words[10]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[10][28] ) );
  DFFX1 \words[10]/data_ff/data_reg[29]  ( .D(\words[10]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[10][29] ) );
  DFFX1 \words[10]/data_ff/data_reg[30]  ( .D(\words[10]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[10][30] ) );
  DFFX1 \words[10]/data_ff/data_reg[31]  ( .D(\words[10]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[10][31] ) );
  DFFX1 \words[11]/data_ff/data_reg[0]  ( .D(\words[11]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[11][0] ) );
  DFFX1 \words[11]/data_ff/data_reg[1]  ( .D(\words[11]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[11][1] ) );
  DFFX1 \words[11]/data_ff/data_reg[2]  ( .D(\words[11]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[11][2] ) );
  DFFX1 \words[11]/data_ff/data_reg[3]  ( .D(\words[11]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[11][3] ) );
  DFFX1 \words[11]/data_ff/data_reg[4]  ( .D(\words[11]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[11][4] ) );
  DFFX1 \words[11]/data_ff/data_reg[5]  ( .D(\words[11]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[11][5] ) );
  DFFX1 \words[11]/data_ff/data_reg[6]  ( .D(\words[11]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[11][6] ) );
  DFFX1 \words[11]/data_ff/data_reg[7]  ( .D(\words[11]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[11][7] ) );
  DFFX1 \words[11]/data_ff/data_reg[8]  ( .D(\words[11]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[11][8] ) );
  DFFX1 \words[11]/data_ff/data_reg[9]  ( .D(\words[11]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[11][9] ) );
  DFFX1 \words[11]/data_ff/data_reg[10]  ( .D(\words[11]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[11][10] ) );
  DFFX1 \words[11]/data_ff/data_reg[11]  ( .D(\words[11]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[11][11] ) );
  DFFX1 \words[11]/data_ff/data_reg[12]  ( .D(\words[11]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[11][12] ) );
  DFFX1 \words[11]/data_ff/data_reg[13]  ( .D(\words[11]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[11][13] ) );
  DFFX1 \words[11]/data_ff/data_reg[14]  ( .D(\words[11]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[11][14] ) );
  DFFX1 \words[11]/data_ff/data_reg[15]  ( .D(\words[11]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[11][15] ) );
  DFFX1 \words[11]/data_ff/data_reg[16]  ( .D(\words[11]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[11][16] ) );
  DFFX1 \words[11]/data_ff/data_reg[17]  ( .D(\words[11]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[11][17] ) );
  DFFX1 \words[11]/data_ff/data_reg[18]  ( .D(\words[11]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[11][18] ) );
  DFFX1 \words[11]/data_ff/data_reg[19]  ( .D(\words[11]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[11][19] ) );
  DFFX1 \words[11]/data_ff/data_reg[20]  ( .D(\words[11]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[11][20] ) );
  DFFX1 \words[11]/data_ff/data_reg[21]  ( .D(\words[11]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[11][21] ) );
  DFFX1 \words[11]/data_ff/data_reg[22]  ( .D(\words[11]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[11][22] ) );
  DFFX1 \words[11]/data_ff/data_reg[23]  ( .D(\words[11]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[11][23] ) );
  DFFX1 \words[11]/data_ff/data_reg[24]  ( .D(\words[11]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[11][24] ) );
  DFFX1 \words[11]/data_ff/data_reg[25]  ( .D(\words[11]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[11][25] ) );
  DFFX1 \words[11]/data_ff/data_reg[26]  ( .D(\words[11]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[11][26] ) );
  DFFX1 \words[11]/data_ff/data_reg[27]  ( .D(\words[11]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[11][27] ) );
  DFFX1 \words[11]/data_ff/data_reg[28]  ( .D(\words[11]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[11][28] ) );
  DFFX1 \words[11]/data_ff/data_reg[29]  ( .D(\words[11]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[11][29] ) );
  DFFX1 \words[11]/data_ff/data_reg[30]  ( .D(\words[11]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[11][30] ) );
  DFFX1 \words[11]/data_ff/data_reg[31]  ( .D(\words[11]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[11][31] ) );
  DFFX1 \words[12]/data_ff/data_reg[0]  ( .D(\words[12]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[12][0] ) );
  DFFX1 \words[12]/data_ff/data_reg[1]  ( .D(\words[12]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[12][1] ) );
  DFFX1 \words[12]/data_ff/data_reg[2]  ( .D(\words[12]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[12][2] ) );
  DFFX1 \words[12]/data_ff/data_reg[3]  ( .D(\words[12]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[12][3] ) );
  DFFX1 \words[12]/data_ff/data_reg[4]  ( .D(\words[12]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[12][4] ) );
  DFFX1 \words[12]/data_ff/data_reg[5]  ( .D(\words[12]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[12][5] ) );
  DFFX1 \words[12]/data_ff/data_reg[6]  ( .D(\words[12]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[12][6] ) );
  DFFX1 \words[12]/data_ff/data_reg[7]  ( .D(\words[12]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[12][7] ) );
  DFFX1 \words[12]/data_ff/data_reg[8]  ( .D(\words[12]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[12][8] ) );
  DFFX1 \words[12]/data_ff/data_reg[9]  ( .D(\words[12]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[12][9] ) );
  DFFX1 \words[12]/data_ff/data_reg[10]  ( .D(\words[12]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[12][10] ) );
  DFFX1 \words[12]/data_ff/data_reg[11]  ( .D(\words[12]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[12][11] ) );
  DFFX1 \words[12]/data_ff/data_reg[12]  ( .D(\words[12]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[12][12] ) );
  DFFX1 \words[12]/data_ff/data_reg[13]  ( .D(\words[12]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[12][13] ) );
  DFFX1 \words[12]/data_ff/data_reg[14]  ( .D(\words[12]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[12][14] ) );
  DFFX1 \words[12]/data_ff/data_reg[15]  ( .D(\words[12]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[12][15] ) );
  DFFX1 \words[12]/data_ff/data_reg[16]  ( .D(\words[12]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[12][16] ) );
  DFFX1 \words[12]/data_ff/data_reg[17]  ( .D(\words[12]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[12][17] ) );
  DFFX1 \words[12]/data_ff/data_reg[18]  ( .D(\words[12]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[12][18] ) );
  DFFX1 \words[12]/data_ff/data_reg[19]  ( .D(\words[12]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[12][19] ) );
  DFFX1 \words[12]/data_ff/data_reg[20]  ( .D(\words[12]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[12][20] ) );
  DFFX1 \words[12]/data_ff/data_reg[21]  ( .D(\words[12]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[12][21] ) );
  DFFX1 \words[12]/data_ff/data_reg[22]  ( .D(\words[12]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[12][22] ) );
  DFFX1 \words[12]/data_ff/data_reg[23]  ( .D(\words[12]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[12][23] ) );
  DFFX1 \words[12]/data_ff/data_reg[24]  ( .D(\words[12]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[12][24] ) );
  DFFX1 \words[12]/data_ff/data_reg[25]  ( .D(\words[12]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[12][25] ) );
  DFFX1 \words[12]/data_ff/data_reg[26]  ( .D(\words[12]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[12][26] ) );
  DFFX1 \words[12]/data_ff/data_reg[27]  ( .D(\words[12]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[12][27] ) );
  DFFX1 \words[12]/data_ff/data_reg[28]  ( .D(\words[12]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[12][28] ) );
  DFFX1 \words[12]/data_ff/data_reg[29]  ( .D(\words[12]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[12][29] ) );
  DFFX1 \words[12]/data_ff/data_reg[30]  ( .D(\words[12]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[12][30] ) );
  DFFX1 \words[12]/data_ff/data_reg[31]  ( .D(\words[12]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[12][31] ) );
  DFFX1 \words[13]/data_ff/data_reg[0]  ( .D(\words[13]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[13][0] ) );
  DFFX1 \words[13]/data_ff/data_reg[1]  ( .D(\words[13]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[13][1] ) );
  DFFX1 \words[13]/data_ff/data_reg[2]  ( .D(\words[13]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[13][2] ) );
  DFFX1 \words[13]/data_ff/data_reg[3]  ( .D(\words[13]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[13][3] ) );
  DFFX1 \words[13]/data_ff/data_reg[4]  ( .D(\words[13]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[13][4] ) );
  DFFX1 \words[13]/data_ff/data_reg[5]  ( .D(\words[13]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[13][5] ) );
  DFFX1 \words[13]/data_ff/data_reg[6]  ( .D(\words[13]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[13][6] ) );
  DFFX1 \words[13]/data_ff/data_reg[7]  ( .D(\words[13]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[13][7] ) );
  DFFX1 \words[13]/data_ff/data_reg[8]  ( .D(\words[13]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[13][8] ) );
  DFFX1 \words[13]/data_ff/data_reg[9]  ( .D(\words[13]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[13][9] ) );
  DFFX1 \words[13]/data_ff/data_reg[10]  ( .D(\words[13]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[13][10] ) );
  DFFX1 \words[13]/data_ff/data_reg[11]  ( .D(\words[13]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[13][11] ) );
  DFFX1 \words[13]/data_ff/data_reg[12]  ( .D(\words[13]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[13][12] ) );
  DFFX1 \words[13]/data_ff/data_reg[13]  ( .D(\words[13]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[13][13] ) );
  DFFX1 \words[13]/data_ff/data_reg[14]  ( .D(\words[13]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[13][14] ) );
  DFFX1 \words[13]/data_ff/data_reg[15]  ( .D(\words[13]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[13][15] ) );
  DFFX1 \words[13]/data_ff/data_reg[16]  ( .D(\words[13]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[13][16] ) );
  DFFX1 \words[13]/data_ff/data_reg[17]  ( .D(\words[13]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[13][17] ) );
  DFFX1 \words[13]/data_ff/data_reg[18]  ( .D(\words[13]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[13][18] ) );
  DFFX1 \words[13]/data_ff/data_reg[19]  ( .D(\words[13]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[13][19] ) );
  DFFX1 \words[13]/data_ff/data_reg[20]  ( .D(\words[13]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[13][20] ) );
  DFFX1 \words[13]/data_ff/data_reg[21]  ( .D(\words[13]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[13][21] ) );
  DFFX1 \words[13]/data_ff/data_reg[22]  ( .D(\words[13]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[13][22] ) );
  DFFX1 \words[13]/data_ff/data_reg[23]  ( .D(\words[13]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[13][23] ) );
  DFFX1 \words[13]/data_ff/data_reg[24]  ( .D(\words[13]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[13][24] ) );
  DFFX1 \words[13]/data_ff/data_reg[25]  ( .D(\words[13]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[13][25] ) );
  DFFX1 \words[13]/data_ff/data_reg[26]  ( .D(\words[13]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[13][26] ) );
  DFFX1 \words[13]/data_ff/data_reg[27]  ( .D(\words[13]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[13][27] ) );
  DFFX1 \words[13]/data_ff/data_reg[28]  ( .D(\words[13]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[13][28] ) );
  DFFX1 \words[13]/data_ff/data_reg[29]  ( .D(\words[13]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[13][29] ) );
  DFFX1 \words[13]/data_ff/data_reg[30]  ( .D(\words[13]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[13][30] ) );
  DFFX1 \words[13]/data_ff/data_reg[31]  ( .D(\words[13]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[13][31] ) );
  DFFX1 \words[14]/data_ff/data_reg[0]  ( .D(\words[14]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[14][0] ) );
  DFFX1 \words[14]/data_ff/data_reg[1]  ( .D(\words[14]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[14][1] ) );
  DFFX1 \words[14]/data_ff/data_reg[2]  ( .D(\words[14]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[14][2] ) );
  DFFX1 \words[14]/data_ff/data_reg[3]  ( .D(\words[14]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[14][3] ) );
  DFFX1 \words[14]/data_ff/data_reg[4]  ( .D(\words[14]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[14][4] ) );
  DFFX1 \words[14]/data_ff/data_reg[5]  ( .D(\words[14]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[14][5] ) );
  DFFX1 \words[14]/data_ff/data_reg[6]  ( .D(\words[14]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[14][6] ) );
  DFFX1 \words[14]/data_ff/data_reg[7]  ( .D(\words[14]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[14][7] ) );
  DFFX1 \words[14]/data_ff/data_reg[8]  ( .D(\words[14]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[14][8] ) );
  DFFX1 \words[14]/data_ff/data_reg[9]  ( .D(\words[14]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[14][9] ) );
  DFFX1 \words[14]/data_ff/data_reg[10]  ( .D(\words[14]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[14][10] ) );
  DFFX1 \words[14]/data_ff/data_reg[11]  ( .D(\words[14]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[14][11] ) );
  DFFX1 \words[14]/data_ff/data_reg[12]  ( .D(\words[14]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[14][12] ) );
  DFFX1 \words[14]/data_ff/data_reg[13]  ( .D(\words[14]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[14][13] ) );
  DFFX1 \words[14]/data_ff/data_reg[14]  ( .D(\words[14]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[14][14] ) );
  DFFX1 \words[14]/data_ff/data_reg[15]  ( .D(\words[14]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[14][15] ) );
  DFFX1 \words[14]/data_ff/data_reg[16]  ( .D(\words[14]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[14][16] ) );
  DFFX1 \words[14]/data_ff/data_reg[17]  ( .D(\words[14]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[14][17] ) );
  DFFX1 \words[14]/data_ff/data_reg[18]  ( .D(\words[14]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[14][18] ) );
  DFFX1 \words[14]/data_ff/data_reg[19]  ( .D(\words[14]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[14][19] ) );
  DFFX1 \words[14]/data_ff/data_reg[20]  ( .D(\words[14]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[14][20] ) );
  DFFX1 \words[14]/data_ff/data_reg[21]  ( .D(\words[14]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[14][21] ) );
  DFFX1 \words[14]/data_ff/data_reg[22]  ( .D(\words[14]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[14][22] ) );
  DFFX1 \words[14]/data_ff/data_reg[23]  ( .D(\words[14]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[14][23] ) );
  DFFX1 \words[14]/data_ff/data_reg[24]  ( .D(\words[14]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[14][24] ) );
  DFFX1 \words[14]/data_ff/data_reg[25]  ( .D(\words[14]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[14][25] ) );
  DFFX1 \words[14]/data_ff/data_reg[26]  ( .D(\words[14]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[14][26] ) );
  DFFX1 \words[14]/data_ff/data_reg[27]  ( .D(\words[14]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[14][27] ) );
  DFFX1 \words[14]/data_ff/data_reg[28]  ( .D(\words[14]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[14][28] ) );
  DFFX1 \words[14]/data_ff/data_reg[29]  ( .D(\words[14]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[14][29] ) );
  DFFX1 \words[14]/data_ff/data_reg[30]  ( .D(\words[14]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[14][30] ) );
  DFFX1 \words[14]/data_ff/data_reg[31]  ( .D(\words[14]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[14][31] ) );
  DFFX1 \words[15]/data_ff/data_reg[0]  ( .D(\words[15]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[15][0] ) );
  DFFX1 \words[15]/data_ff/data_reg[1]  ( .D(\words[15]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[15][1] ) );
  DFFX1 \words[15]/data_ff/data_reg[2]  ( .D(\words[15]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[15][2] ) );
  DFFX1 \words[15]/data_ff/data_reg[3]  ( .D(\words[15]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[15][3] ) );
  DFFX1 \words[15]/data_ff/data_reg[4]  ( .D(\words[15]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[15][4] ) );
  DFFX1 \words[15]/data_ff/data_reg[5]  ( .D(\words[15]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[15][5] ) );
  DFFX1 \words[15]/data_ff/data_reg[6]  ( .D(\words[15]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[15][6] ) );
  DFFX1 \words[15]/data_ff/data_reg[7]  ( .D(\words[15]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[15][7] ) );
  DFFX1 \words[15]/data_ff/data_reg[8]  ( .D(\words[15]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[15][8] ) );
  DFFX1 \words[15]/data_ff/data_reg[9]  ( .D(\words[15]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[15][9] ) );
  DFFX1 \words[15]/data_ff/data_reg[10]  ( .D(\words[15]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[15][10] ) );
  DFFX1 \words[15]/data_ff/data_reg[11]  ( .D(\words[15]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[15][11] ) );
  DFFX1 \words[15]/data_ff/data_reg[12]  ( .D(\words[15]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[15][12] ) );
  DFFX1 \words[15]/data_ff/data_reg[13]  ( .D(\words[15]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[15][13] ) );
  DFFX1 \words[15]/data_ff/data_reg[14]  ( .D(\words[15]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[15][14] ) );
  DFFX1 \words[15]/data_ff/data_reg[15]  ( .D(\words[15]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[15][15] ) );
  DFFX1 \words[15]/data_ff/data_reg[16]  ( .D(\words[15]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[15][16] ) );
  DFFX1 \words[15]/data_ff/data_reg[17]  ( .D(\words[15]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[15][17] ) );
  DFFX1 \words[15]/data_ff/data_reg[18]  ( .D(\words[15]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[15][18] ) );
  DFFX1 \words[15]/data_ff/data_reg[19]  ( .D(\words[15]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[15][19] ) );
  DFFX1 \words[15]/data_ff/data_reg[20]  ( .D(\words[15]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[15][20] ) );
  DFFX1 \words[15]/data_ff/data_reg[21]  ( .D(\words[15]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[15][21] ) );
  DFFX1 \words[15]/data_ff/data_reg[22]  ( .D(\words[15]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[15][22] ) );
  DFFX1 \words[15]/data_ff/data_reg[23]  ( .D(\words[15]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[15][23] ) );
  DFFX1 \words[15]/data_ff/data_reg[24]  ( .D(\words[15]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[15][24] ) );
  DFFX1 \words[15]/data_ff/data_reg[25]  ( .D(\words[15]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[15][25] ) );
  DFFX1 \words[15]/data_ff/data_reg[26]  ( .D(\words[15]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[15][26] ) );
  DFFX1 \words[15]/data_ff/data_reg[27]  ( .D(\words[15]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[15][27] ) );
  DFFX1 \words[15]/data_ff/data_reg[28]  ( .D(\words[15]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[15][28] ) );
  DFFX1 \words[15]/data_ff/data_reg[29]  ( .D(\words[15]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[15][29] ) );
  DFFX1 \words[15]/data_ff/data_reg[30]  ( .D(\words[15]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[15][30] ) );
  DFFX1 \words[15]/data_ff/data_reg[31]  ( .D(\words[15]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[15][31] ) );
  DFFX1 \words[16]/data_ff/data_reg[0]  ( .D(\words[16]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[16][0] ) );
  DFFX1 \words[16]/data_ff/data_reg[1]  ( .D(\words[16]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[16][1] ) );
  DFFX1 \words[16]/data_ff/data_reg[2]  ( .D(\words[16]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[16][2] ) );
  DFFX1 \words[16]/data_ff/data_reg[3]  ( .D(\words[16]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[16][3] ) );
  DFFX1 \words[16]/data_ff/data_reg[4]  ( .D(\words[16]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[16][4] ) );
  DFFX1 \words[16]/data_ff/data_reg[5]  ( .D(\words[16]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[16][5] ) );
  DFFX1 \words[16]/data_ff/data_reg[6]  ( .D(\words[16]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[16][6] ) );
  DFFX1 \words[16]/data_ff/data_reg[7]  ( .D(\words[16]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[16][7] ) );
  DFFX1 \words[16]/data_ff/data_reg[8]  ( .D(\words[16]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[16][8] ) );
  DFFX1 \words[16]/data_ff/data_reg[9]  ( .D(\words[16]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[16][9] ) );
  DFFX1 \words[16]/data_ff/data_reg[10]  ( .D(\words[16]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[16][10] ) );
  DFFX1 \words[16]/data_ff/data_reg[11]  ( .D(\words[16]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[16][11] ) );
  DFFX1 \words[16]/data_ff/data_reg[12]  ( .D(\words[16]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[16][12] ) );
  DFFX1 \words[16]/data_ff/data_reg[13]  ( .D(\words[16]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[16][13] ) );
  DFFX1 \words[16]/data_ff/data_reg[14]  ( .D(\words[16]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[16][14] ) );
  DFFX1 \words[16]/data_ff/data_reg[15]  ( .D(\words[16]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[16][15] ) );
  DFFX1 \words[16]/data_ff/data_reg[16]  ( .D(\words[16]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[16][16] ) );
  DFFX1 \words[16]/data_ff/data_reg[17]  ( .D(\words[16]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[16][17] ) );
  DFFX1 \words[16]/data_ff/data_reg[18]  ( .D(\words[16]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[16][18] ) );
  DFFX1 \words[16]/data_ff/data_reg[19]  ( .D(\words[16]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[16][19] ) );
  DFFX1 \words[16]/data_ff/data_reg[20]  ( .D(\words[16]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[16][20] ) );
  DFFX1 \words[16]/data_ff/data_reg[21]  ( .D(\words[16]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[16][21] ) );
  DFFX1 \words[16]/data_ff/data_reg[22]  ( .D(\words[16]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[16][22] ) );
  DFFX1 \words[16]/data_ff/data_reg[23]  ( .D(\words[16]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[16][23] ) );
  DFFX1 \words[16]/data_ff/data_reg[24]  ( .D(\words[16]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[16][24] ) );
  DFFX1 \words[16]/data_ff/data_reg[25]  ( .D(\words[16]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[16][25] ) );
  DFFX1 \words[16]/data_ff/data_reg[26]  ( .D(\words[16]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[16][26] ) );
  DFFX1 \words[16]/data_ff/data_reg[27]  ( .D(\words[16]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[16][27] ) );
  DFFX1 \words[16]/data_ff/data_reg[28]  ( .D(\words[16]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[16][28] ) );
  DFFX1 \words[16]/data_ff/data_reg[29]  ( .D(\words[16]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[16][29] ) );
  DFFX1 \words[16]/data_ff/data_reg[30]  ( .D(\words[16]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[16][30] ) );
  DFFX1 \words[16]/data_ff/data_reg[31]  ( .D(\words[16]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[16][31] ) );
  DFFX1 \words[17]/data_ff/data_reg[0]  ( .D(\words[17]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[17][0] ) );
  DFFX1 \words[17]/data_ff/data_reg[1]  ( .D(\words[17]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[17][1] ) );
  DFFX1 \words[17]/data_ff/data_reg[2]  ( .D(\words[17]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[17][2] ) );
  DFFX1 \words[17]/data_ff/data_reg[3]  ( .D(\words[17]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[17][3] ) );
  DFFX1 \words[17]/data_ff/data_reg[4]  ( .D(\words[17]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[17][4] ) );
  DFFX1 \words[17]/data_ff/data_reg[5]  ( .D(\words[17]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[17][5] ) );
  DFFX1 \words[17]/data_ff/data_reg[6]  ( .D(\words[17]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[17][6] ) );
  DFFX1 \words[17]/data_ff/data_reg[7]  ( .D(\words[17]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[17][7] ) );
  DFFX1 \words[17]/data_ff/data_reg[8]  ( .D(\words[17]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[17][8] ) );
  DFFX1 \words[17]/data_ff/data_reg[9]  ( .D(\words[17]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[17][9] ) );
  DFFX1 \words[17]/data_ff/data_reg[10]  ( .D(\words[17]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[17][10] ) );
  DFFX1 \words[17]/data_ff/data_reg[11]  ( .D(\words[17]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[17][11] ) );
  DFFX1 \words[17]/data_ff/data_reg[12]  ( .D(\words[17]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[17][12] ) );
  DFFX1 \words[17]/data_ff/data_reg[13]  ( .D(\words[17]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[17][13] ) );
  DFFX1 \words[17]/data_ff/data_reg[14]  ( .D(\words[17]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[17][14] ) );
  DFFX1 \words[17]/data_ff/data_reg[15]  ( .D(\words[17]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[17][15] ) );
  DFFX1 \words[17]/data_ff/data_reg[16]  ( .D(\words[17]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[17][16] ) );
  DFFX1 \words[17]/data_ff/data_reg[17]  ( .D(\words[17]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[17][17] ) );
  DFFX1 \words[17]/data_ff/data_reg[18]  ( .D(\words[17]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[17][18] ) );
  DFFX1 \words[17]/data_ff/data_reg[19]  ( .D(\words[17]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[17][19] ) );
  DFFX1 \words[17]/data_ff/data_reg[20]  ( .D(\words[17]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[17][20] ) );
  DFFX1 \words[17]/data_ff/data_reg[21]  ( .D(\words[17]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[17][21] ) );
  DFFX1 \words[17]/data_ff/data_reg[22]  ( .D(\words[17]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[17][22] ) );
  DFFX1 \words[17]/data_ff/data_reg[23]  ( .D(\words[17]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[17][23] ) );
  DFFX1 \words[17]/data_ff/data_reg[24]  ( .D(\words[17]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[17][24] ) );
  DFFX1 \words[17]/data_ff/data_reg[25]  ( .D(\words[17]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[17][25] ) );
  DFFX1 \words[17]/data_ff/data_reg[26]  ( .D(\words[17]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[17][26] ) );
  DFFX1 \words[17]/data_ff/data_reg[27]  ( .D(\words[17]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[17][27] ) );
  DFFX1 \words[17]/data_ff/data_reg[28]  ( .D(\words[17]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[17][28] ) );
  DFFX1 \words[17]/data_ff/data_reg[29]  ( .D(\words[17]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[17][29] ) );
  DFFX1 \words[17]/data_ff/data_reg[30]  ( .D(\words[17]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[17][30] ) );
  DFFX1 \words[17]/data_ff/data_reg[31]  ( .D(\words[17]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[17][31] ) );
  DFFX1 \words[18]/data_ff/data_reg[0]  ( .D(\words[18]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[18][0] ) );
  DFFX1 \words[18]/data_ff/data_reg[1]  ( .D(\words[18]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[18][1] ) );
  DFFX1 \words[18]/data_ff/data_reg[2]  ( .D(\words[18]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[18][2] ) );
  DFFX1 \words[18]/data_ff/data_reg[3]  ( .D(\words[18]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[18][3] ) );
  DFFX1 \words[18]/data_ff/data_reg[4]  ( .D(\words[18]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[18][4] ) );
  DFFX1 \words[18]/data_ff/data_reg[5]  ( .D(\words[18]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[18][5] ) );
  DFFX1 \words[18]/data_ff/data_reg[6]  ( .D(\words[18]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[18][6] ) );
  DFFX1 \words[18]/data_ff/data_reg[7]  ( .D(\words[18]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[18][7] ) );
  DFFX1 \words[18]/data_ff/data_reg[8]  ( .D(\words[18]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[18][8] ), .QN(n1649) );
  DFFX1 \words[18]/data_ff/data_reg[9]  ( .D(\words[18]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[18][9] ) );
  DFFX1 \words[18]/data_ff/data_reg[10]  ( .D(\words[18]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[18][10] ) );
  DFFX1 \words[18]/data_ff/data_reg[11]  ( .D(\words[18]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[18][11] ) );
  DFFX1 \words[18]/data_ff/data_reg[12]  ( .D(\words[18]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[18][12] ) );
  DFFX1 \words[18]/data_ff/data_reg[13]  ( .D(\words[18]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[18][13] ) );
  DFFX1 \words[18]/data_ff/data_reg[14]  ( .D(\words[18]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[18][14] ) );
  DFFX1 \words[18]/data_ff/data_reg[15]  ( .D(\words[18]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[18][15] ) );
  DFFX1 \words[18]/data_ff/data_reg[16]  ( .D(\words[18]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[18][16] ) );
  DFFX1 \words[18]/data_ff/data_reg[17]  ( .D(\words[18]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[18][17] ) );
  DFFX1 \words[18]/data_ff/data_reg[18]  ( .D(\words[18]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[18][18] ) );
  DFFX1 \words[18]/data_ff/data_reg[19]  ( .D(\words[18]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[18][19] ) );
  DFFX1 \words[18]/data_ff/data_reg[20]  ( .D(\words[18]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[18][20] ) );
  DFFX1 \words[18]/data_ff/data_reg[21]  ( .D(\words[18]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[18][21] ) );
  DFFX1 \words[18]/data_ff/data_reg[22]  ( .D(\words[18]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[18][22] ) );
  DFFX1 \words[18]/data_ff/data_reg[23]  ( .D(\words[18]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[18][23] ) );
  DFFX1 \words[18]/data_ff/data_reg[24]  ( .D(\words[18]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[18][24] ) );
  DFFX1 \words[18]/data_ff/data_reg[25]  ( .D(\words[18]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[18][25] ) );
  DFFX1 \words[18]/data_ff/data_reg[26]  ( .D(\words[18]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[18][26] ) );
  DFFX1 \words[18]/data_ff/data_reg[27]  ( .D(\words[18]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[18][27] ), .QN(n1652) );
  DFFX1 \words[18]/data_ff/data_reg[28]  ( .D(\words[18]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[18][28] ) );
  DFFX1 \words[18]/data_ff/data_reg[29]  ( .D(\words[18]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[18][29] ) );
  DFFX1 \words[18]/data_ff/data_reg[30]  ( .D(\words[18]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[18][30] ) );
  DFFX1 \words[18]/data_ff/data_reg[31]  ( .D(\words[18]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[18][31] ) );
  DFFX1 \words[19]/data_ff/data_reg[0]  ( .D(\words[19]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[19][0] ) );
  DFFX1 \words[19]/data_ff/data_reg[1]  ( .D(\words[19]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[19][1] ) );
  DFFX1 \words[19]/data_ff/data_reg[2]  ( .D(\words[19]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[19][2] ) );
  DFFX1 \words[19]/data_ff/data_reg[3]  ( .D(\words[19]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[19][3] ) );
  DFFX1 \words[19]/data_ff/data_reg[4]  ( .D(\words[19]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[19][4] ) );
  DFFX1 \words[19]/data_ff/data_reg[5]  ( .D(\words[19]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[19][5] ) );
  DFFX1 \words[19]/data_ff/data_reg[6]  ( .D(\words[19]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[19][6] ) );
  DFFX1 \words[19]/data_ff/data_reg[7]  ( .D(\words[19]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[19][7] ) );
  DFFX1 \words[19]/data_ff/data_reg[8]  ( .D(\words[19]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[19][8] ) );
  DFFX1 \words[19]/data_ff/data_reg[9]  ( .D(\words[19]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[19][9] ) );
  DFFX1 \words[19]/data_ff/data_reg[10]  ( .D(\words[19]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[19][10] ) );
  DFFX1 \words[19]/data_ff/data_reg[11]  ( .D(\words[19]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[19][11] ) );
  DFFX1 \words[19]/data_ff/data_reg[12]  ( .D(\words[19]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[19][12] ) );
  DFFX1 \words[19]/data_ff/data_reg[13]  ( .D(\words[19]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[19][13] ) );
  DFFX1 \words[19]/data_ff/data_reg[14]  ( .D(\words[19]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[19][14] ) );
  DFFX1 \words[19]/data_ff/data_reg[15]  ( .D(\words[19]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[19][15] ) );
  DFFX1 \words[19]/data_ff/data_reg[16]  ( .D(\words[19]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[19][16] ) );
  DFFX1 \words[19]/data_ff/data_reg[17]  ( .D(\words[19]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[19][17] ) );
  DFFX1 \words[19]/data_ff/data_reg[18]  ( .D(\words[19]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[19][18] ) );
  DFFX1 \words[19]/data_ff/data_reg[19]  ( .D(\words[19]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[19][19] ) );
  DFFX1 \words[19]/data_ff/data_reg[20]  ( .D(\words[19]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[19][20] ) );
  DFFX1 \words[19]/data_ff/data_reg[21]  ( .D(\words[19]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[19][21] ) );
  DFFX1 \words[19]/data_ff/data_reg[22]  ( .D(\words[19]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[19][22] ) );
  DFFX1 \words[19]/data_ff/data_reg[23]  ( .D(\words[19]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[19][23] ) );
  DFFX1 \words[19]/data_ff/data_reg[24]  ( .D(\words[19]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[19][24] ) );
  DFFX1 \words[19]/data_ff/data_reg[25]  ( .D(\words[19]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[19][25] ) );
  DFFX1 \words[19]/data_ff/data_reg[26]  ( .D(\words[19]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[19][26] ) );
  DFFX1 \words[19]/data_ff/data_reg[27]  ( .D(\words[19]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[19][27] ) );
  DFFX1 \words[19]/data_ff/data_reg[28]  ( .D(\words[19]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[19][28] ) );
  DFFX1 \words[19]/data_ff/data_reg[29]  ( .D(\words[19]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[19][29] ) );
  DFFX1 \words[19]/data_ff/data_reg[30]  ( .D(\words[19]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[19][30] ) );
  DFFX1 \words[19]/data_ff/data_reg[31]  ( .D(\words[19]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[19][31] ) );
  DFFX1 \words[20]/data_ff/data_reg[0]  ( .D(\words[20]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[20][0] ) );
  DFFX1 \words[20]/data_ff/data_reg[1]  ( .D(\words[20]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[20][1] ) );
  DFFX1 \words[20]/data_ff/data_reg[2]  ( .D(\words[20]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[20][2] ) );
  DFFX1 \words[20]/data_ff/data_reg[3]  ( .D(\words[20]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[20][3] ) );
  DFFX1 \words[20]/data_ff/data_reg[4]  ( .D(\words[20]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[20][4] ) );
  DFFX1 \words[20]/data_ff/data_reg[5]  ( .D(\words[20]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[20][5] ) );
  DFFX1 \words[20]/data_ff/data_reg[6]  ( .D(\words[20]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[20][6] ) );
  DFFX1 \words[20]/data_ff/data_reg[7]  ( .D(\words[20]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[20][7] ) );
  DFFX1 \words[20]/data_ff/data_reg[8]  ( .D(\words[20]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[20][8] ) );
  DFFX1 \words[20]/data_ff/data_reg[9]  ( .D(\words[20]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[20][9] ) );
  DFFX1 \words[20]/data_ff/data_reg[10]  ( .D(\words[20]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[20][10] ) );
  DFFX1 \words[20]/data_ff/data_reg[11]  ( .D(\words[20]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[20][11] ) );
  DFFX1 \words[20]/data_ff/data_reg[12]  ( .D(\words[20]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[20][12] ) );
  DFFX1 \words[20]/data_ff/data_reg[13]  ( .D(\words[20]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[20][13] ) );
  DFFX1 \words[20]/data_ff/data_reg[14]  ( .D(\words[20]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[20][14] ) );
  DFFX1 \words[20]/data_ff/data_reg[15]  ( .D(\words[20]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[20][15] ) );
  DFFX1 \words[20]/data_ff/data_reg[16]  ( .D(\words[20]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[20][16] ) );
  DFFX1 \words[20]/data_ff/data_reg[17]  ( .D(\words[20]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[20][17] ) );
  DFFX1 \words[20]/data_ff/data_reg[18]  ( .D(\words[20]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[20][18] ) );
  DFFX1 \words[20]/data_ff/data_reg[19]  ( .D(\words[20]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[20][19] ) );
  DFFX1 \words[20]/data_ff/data_reg[20]  ( .D(\words[20]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[20][20] ) );
  DFFX1 \words[20]/data_ff/data_reg[21]  ( .D(\words[20]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[20][21] ) );
  DFFX1 \words[20]/data_ff/data_reg[22]  ( .D(\words[20]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[20][22] ) );
  DFFX1 \words[20]/data_ff/data_reg[23]  ( .D(\words[20]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[20][23] ) );
  DFFX1 \words[20]/data_ff/data_reg[24]  ( .D(\words[20]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[20][24] ) );
  DFFX1 \words[20]/data_ff/data_reg[25]  ( .D(\words[20]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[20][25] ) );
  DFFX1 \words[20]/data_ff/data_reg[26]  ( .D(\words[20]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[20][26] ) );
  DFFX1 \words[20]/data_ff/data_reg[27]  ( .D(\words[20]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[20][27] ) );
  DFFX1 \words[20]/data_ff/data_reg[28]  ( .D(\words[20]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[20][28] ) );
  DFFX1 \words[20]/data_ff/data_reg[29]  ( .D(\words[20]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[20][29] ) );
  DFFX1 \words[20]/data_ff/data_reg[30]  ( .D(\words[20]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[20][30] ) );
  DFFX1 \words[20]/data_ff/data_reg[31]  ( .D(\words[20]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[20][31] ) );
  DFFX1 \words[21]/data_ff/data_reg[0]  ( .D(\words[21]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[21][0] ) );
  DFFX1 \words[21]/data_ff/data_reg[1]  ( .D(\words[21]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[21][1] ) );
  DFFX1 \words[21]/data_ff/data_reg[2]  ( .D(\words[21]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[21][2] ) );
  DFFX1 \words[21]/data_ff/data_reg[3]  ( .D(\words[21]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[21][3] ) );
  DFFX1 \words[21]/data_ff/data_reg[4]  ( .D(\words[21]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[21][4] ) );
  DFFX1 \words[21]/data_ff/data_reg[5]  ( .D(\words[21]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[21][5] ) );
  DFFX1 \words[21]/data_ff/data_reg[6]  ( .D(\words[21]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[21][6] ) );
  DFFX1 \words[21]/data_ff/data_reg[7]  ( .D(\words[21]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[21][7] ) );
  DFFX1 \words[21]/data_ff/data_reg[8]  ( .D(\words[21]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[21][8] ) );
  DFFX1 \words[21]/data_ff/data_reg[9]  ( .D(\words[21]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[21][9] ) );
  DFFX1 \words[21]/data_ff/data_reg[10]  ( .D(\words[21]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[21][10] ) );
  DFFX1 \words[21]/data_ff/data_reg[11]  ( .D(\words[21]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[21][11] ) );
  DFFX1 \words[21]/data_ff/data_reg[12]  ( .D(\words[21]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[21][12] ) );
  DFFX1 \words[21]/data_ff/data_reg[13]  ( .D(\words[21]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[21][13] ) );
  DFFX1 \words[21]/data_ff/data_reg[14]  ( .D(\words[21]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[21][14] ) );
  DFFX1 \words[21]/data_ff/data_reg[15]  ( .D(\words[21]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[21][15] ) );
  DFFX1 \words[21]/data_ff/data_reg[16]  ( .D(\words[21]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[21][16] ) );
  DFFX1 \words[21]/data_ff/data_reg[17]  ( .D(\words[21]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[21][17] ) );
  DFFX1 \words[21]/data_ff/data_reg[18]  ( .D(\words[21]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[21][18] ) );
  DFFX1 \words[21]/data_ff/data_reg[19]  ( .D(\words[21]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[21][19] ) );
  DFFX1 \words[21]/data_ff/data_reg[20]  ( .D(\words[21]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[21][20] ) );
  DFFX1 \words[21]/data_ff/data_reg[21]  ( .D(\words[21]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[21][21] ) );
  DFFX1 \words[21]/data_ff/data_reg[22]  ( .D(\words[21]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[21][22] ) );
  DFFX1 \words[21]/data_ff/data_reg[23]  ( .D(\words[21]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[21][23] ) );
  DFFX1 \words[21]/data_ff/data_reg[24]  ( .D(\words[21]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[21][24] ) );
  DFFX1 \words[21]/data_ff/data_reg[25]  ( .D(\words[21]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[21][25] ) );
  DFFX1 \words[21]/data_ff/data_reg[26]  ( .D(\words[21]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[21][26] ) );
  DFFX1 \words[21]/data_ff/data_reg[27]  ( .D(\words[21]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[21][27] ) );
  DFFX1 \words[21]/data_ff/data_reg[28]  ( .D(\words[21]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[21][28] ) );
  DFFX1 \words[21]/data_ff/data_reg[29]  ( .D(\words[21]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[21][29] ) );
  DFFX1 \words[21]/data_ff/data_reg[30]  ( .D(\words[21]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[21][30] ) );
  DFFX1 \words[21]/data_ff/data_reg[31]  ( .D(\words[21]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[21][31] ) );
  DFFX1 \words[22]/data_ff/data_reg[0]  ( .D(\words[22]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[22][0] ) );
  DFFX1 \words[22]/data_ff/data_reg[1]  ( .D(\words[22]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[22][1] ) );
  DFFX1 \words[22]/data_ff/data_reg[2]  ( .D(\words[22]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[22][2] ) );
  DFFX1 \words[22]/data_ff/data_reg[3]  ( .D(\words[22]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[22][3] ) );
  DFFX1 \words[22]/data_ff/data_reg[4]  ( .D(\words[22]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[22][4] ) );
  DFFX1 \words[22]/data_ff/data_reg[5]  ( .D(\words[22]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[22][5] ) );
  DFFX1 \words[22]/data_ff/data_reg[6]  ( .D(\words[22]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[22][6] ) );
  DFFX1 \words[22]/data_ff/data_reg[7]  ( .D(\words[22]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[22][7] ) );
  DFFX1 \words[22]/data_ff/data_reg[8]  ( .D(\words[22]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[22][8] ) );
  DFFX1 \words[22]/data_ff/data_reg[9]  ( .D(\words[22]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[22][9] ) );
  DFFX1 \words[22]/data_ff/data_reg[10]  ( .D(\words[22]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[22][10] ) );
  DFFX1 \words[22]/data_ff/data_reg[11]  ( .D(\words[22]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[22][11] ) );
  DFFX1 \words[22]/data_ff/data_reg[12]  ( .D(\words[22]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[22][12] ) );
  DFFX1 \words[22]/data_ff/data_reg[13]  ( .D(\words[22]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[22][13] ) );
  DFFX1 \words[22]/data_ff/data_reg[14]  ( .D(\words[22]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[22][14] ) );
  DFFX1 \words[22]/data_ff/data_reg[15]  ( .D(\words[22]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[22][15] ) );
  DFFX1 \words[22]/data_ff/data_reg[16]  ( .D(\words[22]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[22][16] ) );
  DFFX1 \words[22]/data_ff/data_reg[17]  ( .D(\words[22]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[22][17] ) );
  DFFX1 \words[22]/data_ff/data_reg[18]  ( .D(\words[22]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[22][18] ) );
  DFFX1 \words[22]/data_ff/data_reg[19]  ( .D(\words[22]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[22][19] ) );
  DFFX1 \words[22]/data_ff/data_reg[20]  ( .D(\words[22]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[22][20] ) );
  DFFX1 \words[22]/data_ff/data_reg[21]  ( .D(\words[22]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[22][21] ) );
  DFFX1 \words[22]/data_ff/data_reg[22]  ( .D(\words[22]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[22][22] ) );
  DFFX1 \words[22]/data_ff/data_reg[23]  ( .D(\words[22]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[22][23] ) );
  DFFX1 \words[22]/data_ff/data_reg[24]  ( .D(\words[22]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[22][24] ) );
  DFFX1 \words[22]/data_ff/data_reg[25]  ( .D(\words[22]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[22][25] ) );
  DFFX1 \words[22]/data_ff/data_reg[26]  ( .D(\words[22]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[22][26] ) );
  DFFX1 \words[22]/data_ff/data_reg[27]  ( .D(\words[22]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[22][27] ) );
  DFFX1 \words[22]/data_ff/data_reg[28]  ( .D(\words[22]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[22][28] ) );
  DFFX1 \words[22]/data_ff/data_reg[29]  ( .D(\words[22]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[22][29] ) );
  DFFX1 \words[22]/data_ff/data_reg[30]  ( .D(\words[22]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[22][30] ) );
  DFFX1 \words[22]/data_ff/data_reg[31]  ( .D(\words[22]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[22][31] ) );
  DFFX1 \words[23]/data_ff/data_reg[0]  ( .D(\words[23]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[23][0] ) );
  DFFX1 \words[23]/data_ff/data_reg[1]  ( .D(\words[23]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[23][1] ) );
  DFFX1 \words[23]/data_ff/data_reg[2]  ( .D(\words[23]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[23][2] ) );
  DFFX1 \words[23]/data_ff/data_reg[3]  ( .D(\words[23]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[23][3] ) );
  DFFX1 \words[23]/data_ff/data_reg[4]  ( .D(\words[23]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[23][4] ) );
  DFFX1 \words[23]/data_ff/data_reg[5]  ( .D(\words[23]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[23][5] ) );
  DFFX1 \words[23]/data_ff/data_reg[6]  ( .D(\words[23]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[23][6] ) );
  DFFX1 \words[23]/data_ff/data_reg[7]  ( .D(\words[23]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[23][7] ) );
  DFFX1 \words[23]/data_ff/data_reg[8]  ( .D(\words[23]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[23][8] ) );
  DFFX1 \words[23]/data_ff/data_reg[9]  ( .D(\words[23]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[23][9] ) );
  DFFX1 \words[23]/data_ff/data_reg[10]  ( .D(\words[23]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[23][10] ) );
  DFFX1 \words[23]/data_ff/data_reg[11]  ( .D(\words[23]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[23][11] ) );
  DFFX1 \words[23]/data_ff/data_reg[12]  ( .D(\words[23]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[23][12] ) );
  DFFX1 \words[23]/data_ff/data_reg[13]  ( .D(\words[23]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[23][13] ) );
  DFFX1 \words[23]/data_ff/data_reg[14]  ( .D(\words[23]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[23][14] ) );
  DFFX1 \words[23]/data_ff/data_reg[15]  ( .D(\words[23]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[23][15] ) );
  DFFX1 \words[23]/data_ff/data_reg[16]  ( .D(\words[23]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[23][16] ) );
  DFFX1 \words[23]/data_ff/data_reg[17]  ( .D(\words[23]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[23][17] ) );
  DFFX1 \words[23]/data_ff/data_reg[18]  ( .D(\words[23]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[23][18] ) );
  DFFX1 \words[23]/data_ff/data_reg[19]  ( .D(\words[23]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[23][19] ) );
  DFFX1 \words[23]/data_ff/data_reg[20]  ( .D(\words[23]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[23][20] ) );
  DFFX1 \words[23]/data_ff/data_reg[21]  ( .D(\words[23]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[23][21] ) );
  DFFX1 \words[23]/data_ff/data_reg[22]  ( .D(\words[23]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[23][22] ) );
  DFFX1 \words[23]/data_ff/data_reg[23]  ( .D(\words[23]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[23][23] ) );
  DFFX1 \words[23]/data_ff/data_reg[24]  ( .D(\words[23]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[23][24] ) );
  DFFX1 \words[23]/data_ff/data_reg[25]  ( .D(\words[23]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[23][25] ) );
  DFFX1 \words[23]/data_ff/data_reg[26]  ( .D(\words[23]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[23][26] ) );
  DFFX1 \words[23]/data_ff/data_reg[27]  ( .D(\words[23]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[23][27] ) );
  DFFX1 \words[23]/data_ff/data_reg[28]  ( .D(\words[23]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[23][28] ) );
  DFFX1 \words[23]/data_ff/data_reg[29]  ( .D(\words[23]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[23][29] ) );
  DFFX1 \words[23]/data_ff/data_reg[30]  ( .D(\words[23]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[23][30] ) );
  DFFX1 \words[23]/data_ff/data_reg[31]  ( .D(\words[23]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[23][31] ) );
  DFFX1 \words[24]/data_ff/data_reg[0]  ( .D(\words[24]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[24][0] ) );
  DFFX1 \words[24]/data_ff/data_reg[1]  ( .D(\words[24]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[24][1] ) );
  DFFX1 \words[24]/data_ff/data_reg[2]  ( .D(\words[24]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[24][2] ) );
  DFFX1 \words[24]/data_ff/data_reg[3]  ( .D(\words[24]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[24][3] ) );
  DFFX1 \words[24]/data_ff/data_reg[4]  ( .D(\words[24]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[24][4] ) );
  DFFX1 \words[24]/data_ff/data_reg[5]  ( .D(\words[24]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[24][5] ) );
  DFFX1 \words[24]/data_ff/data_reg[6]  ( .D(\words[24]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[24][6] ) );
  DFFX1 \words[24]/data_ff/data_reg[7]  ( .D(\words[24]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[24][7] ) );
  DFFX1 \words[24]/data_ff/data_reg[8]  ( .D(\words[24]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[24][8] ) );
  DFFX1 \words[24]/data_ff/data_reg[9]  ( .D(\words[24]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[24][9] ) );
  DFFX1 \words[24]/data_ff/data_reg[10]  ( .D(\words[24]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[24][10] ) );
  DFFX1 \words[24]/data_ff/data_reg[11]  ( .D(\words[24]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[24][11] ) );
  DFFX1 \words[24]/data_ff/data_reg[12]  ( .D(\words[24]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[24][12] ) );
  DFFX1 \words[24]/data_ff/data_reg[13]  ( .D(\words[24]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[24][13] ) );
  DFFX1 \words[24]/data_ff/data_reg[14]  ( .D(\words[24]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[24][14] ) );
  DFFX1 \words[24]/data_ff/data_reg[15]  ( .D(\words[24]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[24][15] ) );
  DFFX1 \words[24]/data_ff/data_reg[16]  ( .D(\words[24]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[24][16] ) );
  DFFX1 \words[24]/data_ff/data_reg[17]  ( .D(\words[24]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[24][17] ) );
  DFFX1 \words[24]/data_ff/data_reg[18]  ( .D(\words[24]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[24][18] ) );
  DFFX1 \words[24]/data_ff/data_reg[19]  ( .D(\words[24]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[24][19] ) );
  DFFX1 \words[24]/data_ff/data_reg[20]  ( .D(\words[24]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[24][20] ) );
  DFFX1 \words[24]/data_ff/data_reg[21]  ( .D(\words[24]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[24][21] ) );
  DFFX1 \words[24]/data_ff/data_reg[22]  ( .D(\words[24]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[24][22] ) );
  DFFX1 \words[24]/data_ff/data_reg[23]  ( .D(\words[24]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[24][23] ) );
  DFFX1 \words[24]/data_ff/data_reg[24]  ( .D(\words[24]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[24][24] ) );
  DFFX1 \words[24]/data_ff/data_reg[25]  ( .D(\words[24]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[24][25] ) );
  DFFX1 \words[24]/data_ff/data_reg[26]  ( .D(\words[24]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[24][26] ) );
  DFFX1 \words[24]/data_ff/data_reg[27]  ( .D(\words[24]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[24][27] ) );
  DFFX1 \words[24]/data_ff/data_reg[28]  ( .D(\words[24]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[24][28] ) );
  DFFX1 \words[24]/data_ff/data_reg[29]  ( .D(\words[24]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[24][29] ) );
  DFFX1 \words[24]/data_ff/data_reg[30]  ( .D(\words[24]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[24][30] ) );
  DFFX1 \words[24]/data_ff/data_reg[31]  ( .D(\words[24]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[24][31] ) );
  DFFX1 \words[25]/data_ff/data_reg[0]  ( .D(\words[25]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[25][0] ) );
  DFFX1 \words[25]/data_ff/data_reg[1]  ( .D(\words[25]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[25][1] ) );
  DFFX1 \words[25]/data_ff/data_reg[2]  ( .D(\words[25]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[25][2] ) );
  DFFX1 \words[25]/data_ff/data_reg[3]  ( .D(\words[25]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[25][3] ) );
  DFFX1 \words[25]/data_ff/data_reg[4]  ( .D(\words[25]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[25][4] ) );
  DFFX1 \words[25]/data_ff/data_reg[5]  ( .D(\words[25]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[25][5] ) );
  DFFX1 \words[25]/data_ff/data_reg[6]  ( .D(\words[25]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[25][6] ) );
  DFFX1 \words[25]/data_ff/data_reg[7]  ( .D(\words[25]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[25][7] ) );
  DFFX1 \words[25]/data_ff/data_reg[8]  ( .D(\words[25]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[25][8] ) );
  DFFX1 \words[25]/data_ff/data_reg[9]  ( .D(\words[25]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[25][9] ) );
  DFFX1 \words[25]/data_ff/data_reg[10]  ( .D(\words[25]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[25][10] ) );
  DFFX1 \words[25]/data_ff/data_reg[11]  ( .D(\words[25]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[25][11] ) );
  DFFX1 \words[25]/data_ff/data_reg[12]  ( .D(\words[25]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[25][12] ) );
  DFFX1 \words[25]/data_ff/data_reg[13]  ( .D(\words[25]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[25][13] ) );
  DFFX1 \words[25]/data_ff/data_reg[14]  ( .D(\words[25]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[25][14] ) );
  DFFX1 \words[25]/data_ff/data_reg[15]  ( .D(\words[25]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[25][15] ) );
  DFFX1 \words[25]/data_ff/data_reg[16]  ( .D(\words[25]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[25][16] ) );
  DFFX1 \words[25]/data_ff/data_reg[17]  ( .D(\words[25]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[25][17] ) );
  DFFX1 \words[25]/data_ff/data_reg[18]  ( .D(\words[25]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[25][18] ) );
  DFFX1 \words[25]/data_ff/data_reg[19]  ( .D(\words[25]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[25][19] ) );
  DFFX1 \words[25]/data_ff/data_reg[20]  ( .D(\words[25]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[25][20] ) );
  DFFX1 \words[25]/data_ff/data_reg[21]  ( .D(\words[25]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[25][21] ) );
  DFFX1 \words[25]/data_ff/data_reg[22]  ( .D(\words[25]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[25][22] ) );
  DFFX1 \words[25]/data_ff/data_reg[23]  ( .D(\words[25]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[25][23] ) );
  DFFX1 \words[25]/data_ff/data_reg[24]  ( .D(\words[25]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[25][24] ) );
  DFFX1 \words[25]/data_ff/data_reg[25]  ( .D(\words[25]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[25][25] ) );
  DFFX1 \words[25]/data_ff/data_reg[26]  ( .D(\words[25]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[25][26] ) );
  DFFX1 \words[25]/data_ff/data_reg[27]  ( .D(\words[25]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[25][27] ) );
  DFFX1 \words[25]/data_ff/data_reg[28]  ( .D(\words[25]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[25][28] ) );
  DFFX1 \words[25]/data_ff/data_reg[29]  ( .D(\words[25]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[25][29] ) );
  DFFX1 \words[25]/data_ff/data_reg[30]  ( .D(\words[25]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[25][30] ) );
  DFFX1 \words[25]/data_ff/data_reg[31]  ( .D(\words[25]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[25][31] ) );
  DFFX1 \words[26]/data_ff/data_reg[0]  ( .D(\words[26]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[26][0] ) );
  DFFX1 \words[26]/data_ff/data_reg[1]  ( .D(\words[26]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[26][1] ) );
  DFFX1 \words[26]/data_ff/data_reg[2]  ( .D(\words[26]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[26][2] ) );
  DFFX1 \words[26]/data_ff/data_reg[3]  ( .D(\words[26]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[26][3] ) );
  DFFX1 \words[26]/data_ff/data_reg[4]  ( .D(\words[26]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[26][4] ) );
  DFFX1 \words[26]/data_ff/data_reg[5]  ( .D(\words[26]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[26][5] ) );
  DFFX1 \words[26]/data_ff/data_reg[6]  ( .D(\words[26]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[26][6] ) );
  DFFX1 \words[26]/data_ff/data_reg[7]  ( .D(\words[26]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[26][7] ) );
  DFFX1 \words[26]/data_ff/data_reg[8]  ( .D(\words[26]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[26][8] ) );
  DFFX1 \words[26]/data_ff/data_reg[9]  ( .D(\words[26]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[26][9] ) );
  DFFX1 \words[26]/data_ff/data_reg[10]  ( .D(\words[26]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[26][10] ) );
  DFFX1 \words[26]/data_ff/data_reg[11]  ( .D(\words[26]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[26][11] ) );
  DFFX1 \words[26]/data_ff/data_reg[12]  ( .D(\words[26]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[26][12] ) );
  DFFX1 \words[26]/data_ff/data_reg[13]  ( .D(\words[26]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[26][13] ) );
  DFFX1 \words[26]/data_ff/data_reg[14]  ( .D(\words[26]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[26][14] ) );
  DFFX1 \words[26]/data_ff/data_reg[15]  ( .D(\words[26]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[26][15] ) );
  DFFX1 \words[26]/data_ff/data_reg[16]  ( .D(\words[26]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[26][16] ) );
  DFFX1 \words[26]/data_ff/data_reg[17]  ( .D(\words[26]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[26][17] ) );
  DFFX1 \words[26]/data_ff/data_reg[18]  ( .D(\words[26]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[26][18] ) );
  DFFX1 \words[26]/data_ff/data_reg[19]  ( .D(\words[26]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[26][19] ) );
  DFFX1 \words[26]/data_ff/data_reg[20]  ( .D(\words[26]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[26][20] ) );
  DFFX1 \words[26]/data_ff/data_reg[21]  ( .D(\words[26]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[26][21] ), .QN(n1653) );
  DFFX1 \words[26]/data_ff/data_reg[22]  ( .D(\words[26]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[26][22] ) );
  DFFX1 \words[26]/data_ff/data_reg[23]  ( .D(\words[26]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[26][23] ) );
  DFFX1 \words[26]/data_ff/data_reg[24]  ( .D(\words[26]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[26][24] ) );
  DFFX1 \words[26]/data_ff/data_reg[25]  ( .D(\words[26]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[26][25] ) );
  DFFX1 \words[26]/data_ff/data_reg[26]  ( .D(\words[26]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[26][26] ) );
  DFFX1 \words[26]/data_ff/data_reg[27]  ( .D(\words[26]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[26][27] ) );
  DFFX1 \words[26]/data_ff/data_reg[28]  ( .D(\words[26]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[26][28] ) );
  DFFX1 \words[26]/data_ff/data_reg[29]  ( .D(\words[26]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[26][29] ) );
  DFFX1 \words[26]/data_ff/data_reg[30]  ( .D(\words[26]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[26][30] ) );
  DFFX1 \words[26]/data_ff/data_reg[31]  ( .D(\words[26]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[26][31] ) );
  DFFX1 \words[27]/data_ff/data_reg[0]  ( .D(\words[27]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[27][0] ) );
  DFFX1 \words[27]/data_ff/data_reg[1]  ( .D(\words[27]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[27][1] ) );
  DFFX1 \words[27]/data_ff/data_reg[2]  ( .D(\words[27]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[27][2] ) );
  DFFX1 \words[27]/data_ff/data_reg[3]  ( .D(\words[27]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[27][3] ) );
  DFFX1 \words[27]/data_ff/data_reg[4]  ( .D(\words[27]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[27][4] ) );
  DFFX1 \words[27]/data_ff/data_reg[5]  ( .D(\words[27]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[27][5] ) );
  DFFX1 \words[27]/data_ff/data_reg[6]  ( .D(\words[27]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[27][6] ) );
  DFFX1 \words[27]/data_ff/data_reg[7]  ( .D(\words[27]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[27][7] ) );
  DFFX1 \words[27]/data_ff/data_reg[8]  ( .D(\words[27]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[27][8] ) );
  DFFX1 \words[27]/data_ff/data_reg[9]  ( .D(\words[27]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[27][9] ) );
  DFFX1 \words[27]/data_ff/data_reg[10]  ( .D(\words[27]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[27][10] ) );
  DFFX1 \words[27]/data_ff/data_reg[11]  ( .D(\words[27]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[27][11] ) );
  DFFX1 \words[27]/data_ff/data_reg[12]  ( .D(\words[27]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[27][12] ) );
  DFFX1 \words[27]/data_ff/data_reg[13]  ( .D(\words[27]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[27][13] ) );
  DFFX1 \words[27]/data_ff/data_reg[14]  ( .D(\words[27]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[27][14] ) );
  DFFX1 \words[27]/data_ff/data_reg[15]  ( .D(\words[27]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[27][15] ) );
  DFFX1 \words[27]/data_ff/data_reg[16]  ( .D(\words[27]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[27][16] ) );
  DFFX1 \words[27]/data_ff/data_reg[17]  ( .D(\words[27]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[27][17] ) );
  DFFX1 \words[27]/data_ff/data_reg[18]  ( .D(\words[27]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[27][18] ) );
  DFFX1 \words[27]/data_ff/data_reg[19]  ( .D(\words[27]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[27][19] ) );
  DFFX1 \words[27]/data_ff/data_reg[20]  ( .D(\words[27]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[27][20] ) );
  DFFX1 \words[27]/data_ff/data_reg[21]  ( .D(\words[27]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[27][21] ) );
  DFFX1 \words[27]/data_ff/data_reg[22]  ( .D(\words[27]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[27][22] ) );
  DFFX1 \words[27]/data_ff/data_reg[23]  ( .D(\words[27]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[27][23] ) );
  DFFX1 \words[27]/data_ff/data_reg[24]  ( .D(\words[27]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[27][24] ) );
  DFFX1 \words[27]/data_ff/data_reg[25]  ( .D(\words[27]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[27][25] ) );
  DFFX1 \words[27]/data_ff/data_reg[26]  ( .D(\words[27]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[27][26] ) );
  DFFX1 \words[27]/data_ff/data_reg[27]  ( .D(\words[27]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[27][27] ) );
  DFFX1 \words[27]/data_ff/data_reg[28]  ( .D(\words[27]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[27][28] ) );
  DFFX1 \words[27]/data_ff/data_reg[29]  ( .D(\words[27]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[27][29] ) );
  DFFX1 \words[27]/data_ff/data_reg[30]  ( .D(\words[27]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[27][30] ) );
  DFFX1 \words[27]/data_ff/data_reg[31]  ( .D(\words[27]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[27][31] ) );
  DFFX1 \words[28]/data_ff/data_reg[0]  ( .D(\words[28]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[28][0] ) );
  DFFX1 \words[28]/data_ff/data_reg[1]  ( .D(\words[28]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[28][1] ) );
  DFFX1 \words[28]/data_ff/data_reg[2]  ( .D(\words[28]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[28][2] ) );
  DFFX1 \words[28]/data_ff/data_reg[3]  ( .D(\words[28]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[28][3] ) );
  DFFX1 \words[28]/data_ff/data_reg[4]  ( .D(\words[28]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[28][4] ) );
  DFFX1 \words[28]/data_ff/data_reg[5]  ( .D(\words[28]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[28][5] ) );
  DFFX1 \words[28]/data_ff/data_reg[6]  ( .D(\words[28]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[28][6] ) );
  DFFX1 \words[28]/data_ff/data_reg[7]  ( .D(\words[28]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[28][7] ) );
  DFFX1 \words[28]/data_ff/data_reg[8]  ( .D(\words[28]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[28][8] ) );
  DFFX1 \words[28]/data_ff/data_reg[9]  ( .D(\words[28]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[28][9] ) );
  DFFX1 \words[28]/data_ff/data_reg[10]  ( .D(\words[28]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[28][10] ) );
  DFFX1 \words[28]/data_ff/data_reg[11]  ( .D(\words[28]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[28][11] ) );
  DFFX1 \words[28]/data_ff/data_reg[12]  ( .D(\words[28]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[28][12] ) );
  DFFX1 \words[28]/data_ff/data_reg[13]  ( .D(\words[28]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[28][13] ) );
  DFFX1 \words[28]/data_ff/data_reg[14]  ( .D(\words[28]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[28][14] ) );
  DFFX1 \words[28]/data_ff/data_reg[15]  ( .D(\words[28]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[28][15] ) );
  DFFX1 \words[28]/data_ff/data_reg[16]  ( .D(\words[28]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[28][16] ) );
  DFFX1 \words[28]/data_ff/data_reg[17]  ( .D(\words[28]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[28][17] ) );
  DFFX1 \words[28]/data_ff/data_reg[18]  ( .D(\words[28]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[28][18] ) );
  DFFX1 \words[28]/data_ff/data_reg[19]  ( .D(\words[28]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[28][19] ) );
  DFFX1 \words[28]/data_ff/data_reg[20]  ( .D(\words[28]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[28][20] ) );
  DFFX1 \words[28]/data_ff/data_reg[21]  ( .D(\words[28]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[28][21] ) );
  DFFX1 \words[28]/data_ff/data_reg[22]  ( .D(\words[28]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[28][22] ) );
  DFFX1 \words[28]/data_ff/data_reg[23]  ( .D(\words[28]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[28][23] ) );
  DFFX1 \words[28]/data_ff/data_reg[24]  ( .D(\words[28]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[28][24] ) );
  DFFX1 \words[28]/data_ff/data_reg[25]  ( .D(\words[28]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[28][25] ) );
  DFFX1 \words[28]/data_ff/data_reg[26]  ( .D(\words[28]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[28][26] ) );
  DFFX1 \words[28]/data_ff/data_reg[27]  ( .D(\words[28]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[28][27] ) );
  DFFX1 \words[28]/data_ff/data_reg[28]  ( .D(\words[28]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[28][28] ) );
  DFFX1 \words[28]/data_ff/data_reg[29]  ( .D(\words[28]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[28][29] ) );
  DFFX1 \words[28]/data_ff/data_reg[30]  ( .D(\words[28]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[28][30] ) );
  DFFX1 \words[28]/data_ff/data_reg[31]  ( .D(\words[28]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[28][31] ) );
  DFFX1 \words[29]/data_ff/data_reg[0]  ( .D(\words[29]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[29][0] ) );
  DFFX1 \words[29]/data_ff/data_reg[1]  ( .D(\words[29]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[29][1] ) );
  DFFX1 \words[29]/data_ff/data_reg[2]  ( .D(\words[29]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[29][2] ) );
  DFFX1 \words[29]/data_ff/data_reg[3]  ( .D(\words[29]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[29][3] ) );
  DFFX1 \words[29]/data_ff/data_reg[4]  ( .D(\words[29]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[29][4] ) );
  DFFX1 \words[29]/data_ff/data_reg[5]  ( .D(\words[29]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[29][5] ) );
  DFFX1 \words[29]/data_ff/data_reg[6]  ( .D(\words[29]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[29][6] ) );
  DFFX1 \words[29]/data_ff/data_reg[7]  ( .D(\words[29]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[29][7] ) );
  DFFX1 \words[29]/data_ff/data_reg[8]  ( .D(\words[29]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[29][8] ) );
  DFFX1 \words[29]/data_ff/data_reg[9]  ( .D(\words[29]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[29][9] ) );
  DFFX1 \words[29]/data_ff/data_reg[10]  ( .D(\words[29]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[29][10] ) );
  DFFX1 \words[29]/data_ff/data_reg[11]  ( .D(\words[29]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[29][11] ) );
  DFFX1 \words[29]/data_ff/data_reg[12]  ( .D(\words[29]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[29][12] ) );
  DFFX1 \words[29]/data_ff/data_reg[13]  ( .D(\words[29]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[29][13] ) );
  DFFX1 \words[29]/data_ff/data_reg[14]  ( .D(\words[29]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[29][14] ) );
  DFFX1 \words[29]/data_ff/data_reg[15]  ( .D(\words[29]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[29][15] ) );
  DFFX1 \words[29]/data_ff/data_reg[16]  ( .D(\words[29]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[29][16] ) );
  DFFX1 \words[29]/data_ff/data_reg[17]  ( .D(\words[29]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[29][17] ) );
  DFFX1 \words[29]/data_ff/data_reg[18]  ( .D(\words[29]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[29][18] ) );
  DFFX1 \words[29]/data_ff/data_reg[19]  ( .D(\words[29]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[29][19] ) );
  DFFX1 \words[29]/data_ff/data_reg[20]  ( .D(\words[29]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[29][20] ) );
  DFFX1 \words[29]/data_ff/data_reg[21]  ( .D(\words[29]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[29][21] ) );
  DFFX1 \words[29]/data_ff/data_reg[22]  ( .D(\words[29]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[29][22] ) );
  DFFX1 \words[29]/data_ff/data_reg[23]  ( .D(\words[29]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[29][23] ) );
  DFFX1 \words[29]/data_ff/data_reg[24]  ( .D(\words[29]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[29][24] ) );
  DFFX1 \words[29]/data_ff/data_reg[25]  ( .D(\words[29]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[29][25] ) );
  DFFX1 \words[29]/data_ff/data_reg[26]  ( .D(\words[29]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[29][26] ) );
  DFFX1 \words[29]/data_ff/data_reg[27]  ( .D(\words[29]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[29][27] ) );
  DFFX1 \words[29]/data_ff/data_reg[28]  ( .D(\words[29]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[29][28] ) );
  DFFX1 \words[29]/data_ff/data_reg[29]  ( .D(\words[29]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[29][29] ) );
  DFFX1 \words[29]/data_ff/data_reg[30]  ( .D(\words[29]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[29][30] ) );
  DFFX1 \words[29]/data_ff/data_reg[31]  ( .D(\words[29]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[29][31] ) );
  DFFX1 \words[30]/data_ff/data_reg[0]  ( .D(\words[30]/data_i[0] ), .CLK(clk), 
        .Q(\read_value_mux[30][0] ) );
  DFFX1 \words[30]/data_ff/data_reg[1]  ( .D(\words[30]/data_i[1] ), .CLK(clk), 
        .Q(\read_value_mux[30][1] ) );
  DFFX1 \words[30]/data_ff/data_reg[2]  ( .D(\words[30]/data_i[2] ), .CLK(clk), 
        .Q(\read_value_mux[30][2] ) );
  DFFX1 \words[30]/data_ff/data_reg[3]  ( .D(\words[30]/data_i[3] ), .CLK(clk), 
        .Q(\read_value_mux[30][3] ) );
  DFFX1 \words[30]/data_ff/data_reg[4]  ( .D(\words[30]/data_i[4] ), .CLK(clk), 
        .Q(\read_value_mux[30][4] ) );
  DFFX1 \words[30]/data_ff/data_reg[5]  ( .D(\words[30]/data_i[5] ), .CLK(clk), 
        .Q(\read_value_mux[30][5] ) );
  DFFX1 \words[30]/data_ff/data_reg[6]  ( .D(\words[30]/data_i[6] ), .CLK(clk), 
        .Q(\read_value_mux[30][6] ) );
  DFFX1 \words[30]/data_ff/data_reg[7]  ( .D(\words[30]/data_i[7] ), .CLK(clk), 
        .Q(\read_value_mux[30][7] ) );
  DFFX1 \words[30]/data_ff/data_reg[8]  ( .D(\words[30]/data_i[8] ), .CLK(clk), 
        .Q(\read_value_mux[30][8] ) );
  DFFX1 \words[30]/data_ff/data_reg[9]  ( .D(\words[30]/data_i[9] ), .CLK(clk), 
        .Q(\read_value_mux[30][9] ) );
  DFFX1 \words[30]/data_ff/data_reg[10]  ( .D(\words[30]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[30][10] ) );
  DFFX1 \words[30]/data_ff/data_reg[11]  ( .D(\words[30]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[30][11] ) );
  DFFX1 \words[30]/data_ff/data_reg[12]  ( .D(\words[30]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[30][12] ) );
  DFFX1 \words[30]/data_ff/data_reg[13]  ( .D(\words[30]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[30][13] ) );
  DFFX1 \words[30]/data_ff/data_reg[14]  ( .D(\words[30]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[30][14] ) );
  DFFX1 \words[30]/data_ff/data_reg[15]  ( .D(\words[30]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[30][15] ) );
  DFFX1 \words[30]/data_ff/data_reg[16]  ( .D(\words[30]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[30][16] ) );
  DFFX1 \words[30]/data_ff/data_reg[17]  ( .D(\words[30]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[30][17] ) );
  DFFX1 \words[30]/data_ff/data_reg[18]  ( .D(\words[30]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[30][18] ) );
  DFFX1 \words[30]/data_ff/data_reg[19]  ( .D(\words[30]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[30][19] ) );
  DFFX1 \words[30]/data_ff/data_reg[20]  ( .D(\words[30]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[30][20] ) );
  DFFX1 \words[30]/data_ff/data_reg[21]  ( .D(\words[30]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[30][21] ) );
  DFFX1 \words[30]/data_ff/data_reg[22]  ( .D(\words[30]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[30][22] ) );
  DFFX1 \words[30]/data_ff/data_reg[23]  ( .D(\words[30]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[30][23] ) );
  DFFX1 \words[30]/data_ff/data_reg[24]  ( .D(\words[30]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[30][24] ) );
  DFFX1 \words[30]/data_ff/data_reg[25]  ( .D(\words[30]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[30][25] ) );
  DFFX1 \words[30]/data_ff/data_reg[26]  ( .D(\words[30]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[30][26] ) );
  DFFX1 \words[30]/data_ff/data_reg[27]  ( .D(\words[30]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[30][27] ) );
  DFFX1 \words[30]/data_ff/data_reg[28]  ( .D(\words[30]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[30][28] ) );
  DFFX1 \words[30]/data_ff/data_reg[29]  ( .D(\words[30]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[30][29] ) );
  DFFX1 \words[30]/data_ff/data_reg[30]  ( .D(\words[30]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[30][30] ) );
  DFFX1 \words[30]/data_ff/data_reg[31]  ( .D(\words[30]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[30][31] ) );
  DFFX1 \words[0]/valid_ff/data_reg[0]  ( .D(\words[0]/valid_i ), .CLK(clk), 
        .Q(\words[0]/valid_o ) );
  DFFX1 \words[1]/valid_ff/data_reg[0]  ( .D(\words[1]/valid_i ), .CLK(clk), 
        .Q(\words[1]/valid_o ) );
  DFFX1 \words[2]/valid_ff/data_reg[0]  ( .D(\words[2]/valid_i ), .CLK(clk), 
        .Q(\words[2]/valid_o ) );
  DFFX1 \words[3]/valid_ff/data_reg[0]  ( .D(\words[3]/valid_i ), .CLK(clk), 
        .Q(\words[3]/valid_o ) );
  DFFX1 \words[4]/valid_ff/data_reg[0]  ( .D(\words[4]/valid_i ), .CLK(clk), 
        .Q(\words[4]/valid_o ) );
  DFFX1 \words[5]/valid_ff/data_reg[0]  ( .D(\words[5]/valid_i ), .CLK(clk), 
        .Q(\words[5]/valid_o ) );
  DFFX1 \words[6]/valid_ff/data_reg[0]  ( .D(\words[6]/valid_i ), .CLK(clk), 
        .Q(\words[6]/valid_o ) );
  DFFX1 \words[7]/valid_ff/data_reg[0]  ( .D(\words[7]/valid_i ), .CLK(clk), 
        .Q(\words[7]/valid_o ) );
  DFFX1 \words[8]/valid_ff/data_reg[0]  ( .D(\words[8]/valid_i ), .CLK(clk), 
        .Q(\words[8]/valid_o ) );
  DFFX1 \words[9]/valid_ff/data_reg[0]  ( .D(\words[9]/valid_i ), .CLK(clk), 
        .Q(\words[9]/valid_o ) );
  DFFX1 \words[10]/valid_ff/data_reg[0]  ( .D(\words[10]/valid_i ), .CLK(clk), 
        .Q(\words[10]/valid_o ) );
  DFFX1 \words[11]/valid_ff/data_reg[0]  ( .D(\words[11]/valid_i ), .CLK(clk), 
        .Q(\words[11]/valid_o ) );
  DFFX1 \words[12]/valid_ff/data_reg[0]  ( .D(\words[12]/valid_i ), .CLK(clk), 
        .Q(\words[12]/valid_o ) );
  DFFX1 \words[13]/valid_ff/data_reg[0]  ( .D(\words[13]/valid_i ), .CLK(clk), 
        .Q(\words[13]/valid_o ) );
  DFFX1 \words[14]/valid_ff/data_reg[0]  ( .D(\words[14]/valid_i ), .CLK(clk), 
        .Q(\words[14]/valid_o ) );
  DFFX1 \words[15]/valid_ff/data_reg[0]  ( .D(\words[15]/valid_i ), .CLK(clk), 
        .Q(\words[15]/valid_o ) );
  DFFX1 \words[16]/valid_ff/data_reg[0]  ( .D(\words[16]/valid_i ), .CLK(clk), 
        .Q(\words[16]/valid_o ) );
  DFFX1 \words[17]/valid_ff/data_reg[0]  ( .D(\words[17]/valid_i ), .CLK(clk), 
        .Q(\words[17]/valid_o ) );
  DFFX1 \words[18]/valid_ff/data_reg[0]  ( .D(\words[18]/valid_i ), .CLK(clk), 
        .Q(\words[18]/valid_o ) );
  DFFX1 \words[19]/valid_ff/data_reg[0]  ( .D(\words[19]/valid_i ), .CLK(clk), 
        .Q(\words[19]/valid_o ) );
  DFFX1 \words[20]/valid_ff/data_reg[0]  ( .D(\words[20]/valid_i ), .CLK(clk), 
        .Q(\words[20]/valid_o ) );
  DFFX1 \words[21]/valid_ff/data_reg[0]  ( .D(\words[21]/valid_i ), .CLK(clk), 
        .Q(\words[21]/valid_o ) );
  DFFX1 \words[22]/valid_ff/data_reg[0]  ( .D(\words[22]/valid_i ), .CLK(clk), 
        .Q(\words[22]/valid_o ) );
  DFFX1 \words[23]/valid_ff/data_reg[0]  ( .D(\words[23]/valid_i ), .CLK(clk), 
        .Q(\words[23]/valid_o ) );
  DFFX1 \words[24]/valid_ff/data_reg[0]  ( .D(\words[24]/valid_i ), .CLK(clk), 
        .Q(\words[24]/valid_o ) );
  DFFX1 \words[25]/valid_ff/data_reg[0]  ( .D(\words[25]/valid_i ), .CLK(clk), 
        .Q(\words[25]/valid_o ) );
  DFFX1 \words[26]/valid_ff/data_reg[0]  ( .D(\words[26]/valid_i ), .CLK(clk), 
        .Q(\words[26]/valid_o ) );
  DFFX1 \words[27]/valid_ff/data_reg[0]  ( .D(\words[27]/valid_i ), .CLK(clk), 
        .Q(\words[27]/valid_o ) );
  DFFX1 \words[28]/valid_ff/data_reg[0]  ( .D(\words[28]/valid_i ), .CLK(clk), 
        .Q(\words[28]/valid_o ) );
  DFFX1 \words[29]/valid_ff/data_reg[0]  ( .D(\words[29]/valid_i ), .CLK(clk), 
        .Q(\words[29]/valid_o ) );
  DFFX1 \words[30]/valid_ff/data_reg[0]  ( .D(\words[30]/valid_i ), .CLK(clk), 
        .Q(\words[30]/valid_o ) );
  MUX21X1 U2646 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[23][28] ), .Q(n2402) );
  MUX21X1 U2647 ( .IN1(n1718), .IN2(search_data[20]), .S(
        \read_value_mux[31][20] ), .Q(n2619) );
  MUX21X1 U2648 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[21][28] ), .Q(n2368) );
  MUX21X1 U2649 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[18][28] ), .Q(n2277) );
  MUX21X1 U2650 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[20][28] ), .Q(n2316) );
  MUX21X1 U2651 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[9][28] ), .Q(n2097) );
  MUX21X1 U2652 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[8][28] ), .Q(n3032) );
  MUX21X1 U2653 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[4][28] ), .Q(n2007) );
  MUX21X1 U2654 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[0][28] ), .Q(n1758) );
  MUX21X1 U2655 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[2][28] ), .Q(n1814) );
  INVX0 U2656 ( .INP(search_data[10]), .ZN(n1691) );
  NOR4X0 U2657 ( .IN1(n2630), .IN2(n2633), .IN3(n2631), .IN4(n2632), .QN(n3074) );
  MUX21X1 U2658 ( .IN1(search_data[31]), .IN2(n1740), .S(
        \read_value_mux[3][31] ), .Q(n1583) );
  MUX21X1 U2659 ( .IN1(search_data[14]), .IN2(n1701), .S(
        \read_value_mux[3][14] ), .Q(n1584) );
  MUX21X1 U2660 ( .IN1(n1676), .IN2(search_data[5]), .S(\read_value_mux[3][5] ), .Q(n1585) );
  MUX21X1 U2661 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[3][28] ), .Q(n1586) );
  MUX21X1 U2662 ( .IN1(n1700), .IN2(search_data[13]), .S(
        \read_value_mux[3][13] ), .Q(n1587) );
  MUX21X1 U2663 ( .IN1(n1716), .IN2(search_data[19]), .S(
        \read_value_mux[3][19] ), .Q(n1588) );
  NAND4X0 U2664 ( .IN1(n1585), .IN2(n1586), .IN3(n1587), .IN4(n1588), .QN(
        n1589) );
  NOR4X0 U2665 ( .IN1(n1659), .IN2(n1583), .IN3(n1584), .IN4(n1589), .QN(n1866) );
  MUX21X1 U2666 ( .IN1(search_data[0]), .IN2(n1661), .S(
        \read_value_mux[29][0] ), .Q(n1590) );
  MUX21X1 U2667 ( .IN1(n1690), .IN2(n1691), .S(\read_value_mux[29][10] ), .Q(
        n1591) );
  MUX21X1 U2668 ( .IN1(n1722), .IN2(search_data[22]), .S(
        \read_value_mux[29][22] ), .Q(n1592) );
  MUX21X1 U2669 ( .IN1(n1682), .IN2(search_data[7]), .S(
        \read_value_mux[29][7] ), .Q(n1593) );
  NAND4X0 U2670 ( .IN1(n1592), .IN2(n2566), .IN3(n1593), .IN4(n2567), .QN(
        n1594) );
  NOR4X0 U2671 ( .IN1(n1611), .IN2(n1590), .IN3(n1591), .IN4(n1594), .QN(n2591) );
  MUX21X1 U2672 ( .IN1(search_data[26]), .IN2(n1728), .S(
        \read_value_mux[25][26] ), .Q(n1595) );
  MUX21X1 U2673 ( .IN1(search_data[25]), .IN2(n1727), .S(
        \read_value_mux[25][25] ), .Q(n1596) );
  NOR4X0 U2674 ( .IN1(n2754), .IN2(n2753), .IN3(n1595), .IN4(n1596), .QN(n3080) );
  MUX21X1 U2675 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[7][28] ), .Q(n1597) );
  MUX21X1 U2676 ( .IN1(n1741), .IN2(search_data[31]), .S(
        \read_value_mux[7][31] ), .Q(n1598) );
  MUX21X1 U2677 ( .IN1(n1696), .IN2(search_data[12]), .S(
        \read_value_mux[7][12] ), .Q(n1599) );
  MUX21X1 U2678 ( .IN1(n1694), .IN2(search_data[11]), .S(
        \read_value_mux[7][11] ), .Q(n1600) );
  NAND4X0 U2679 ( .IN1(n1597), .IN2(n1598), .IN3(n1599), .IN4(n1600), .QN(
        n1938) );
  MUX21X1 U2680 ( .IN1(n1676), .IN2(search_data[5]), .S(
        \read_value_mux[12][5] ), .Q(n1601) );
  MUX21X1 U2681 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[12][25] ), .Q(n1602) );
  MUX21X1 U2682 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[12][28] ), .Q(n1603) );
  MUX21X1 U2683 ( .IN1(n1710), .IN2(search_data[17]), .S(
        \read_value_mux[12][17] ), .Q(n1604) );
  NAND4X0 U2684 ( .IN1(n1601), .IN2(n1602), .IN3(n1603), .IN4(n1604), .QN(
        n2237) );
  INVX0 U2685 ( .INP(n1612), .ZN(n1605) );
  NOR2X0 U2686 ( .IN1(n3109), .IN2(n1605), .QN(n3130) );
  NAND4X0 U2687 ( .IN1(n2562), .IN2(n2563), .IN3(n2564), .IN4(n2565), .QN(
        n1606) );
  NAND3X0 U2688 ( .IN1(n2590), .IN2(n2591), .IN3(n1613), .QN(n1607) );
  NOR4X0 U2689 ( .IN1(n2593), .IN2(n2592), .IN3(n1606), .IN4(n1607), .QN(n3077) );
  OA221X1 U2690 ( .IN1(n3058), .IN2(n3060), .IN3(n3058), .IN4(n3061), .IN5(
        n3057), .Q(n1608) );
  AO221X1 U2691 ( .IN1(n3013), .IN2(n3117), .IN3(n3013), .IN4(n1608), .IN5(
        n3118), .Q(n1609) );
  AO22X1 U2692 ( .IN1(n1654), .IN2(n1655), .IN3(n3056), .IN4(n1609), .Q(
        search_index[0]) );
  INVX0 U2693 ( .INP(n3139), .ZN(n1610) );
  NAND3X0 U2694 ( .IN1(n3140), .IN2(n3138), .IN3(n1610), .QN(search_valid) );
  IBUFFX4 U2695 ( .INP(search_data[20]), .ZN(n1718) );
  NOR2X1 U2696 ( .IN1(reset), .IN2(n3143), .QN(n1623) );
  NOR2X1 U2697 ( .IN1(reset), .IN2(n3165), .QN(n1630) );
  NOR2X1 U2698 ( .IN1(reset), .IN2(n3166), .QN(n1631) );
  NOR2X1 U2699 ( .IN1(reset), .IN2(n3167), .QN(n1639) );
  NOR2X1 U2700 ( .IN1(reset), .IN2(n3169), .QN(n1640) );
  NOR2X1 U2701 ( .IN1(reset), .IN2(n3171), .QN(n1632) );
  NOR2X1 U2702 ( .IN1(reset), .IN2(n3172), .QN(n1633) );
  NOR2X1 U2703 ( .IN1(reset), .IN2(n3174), .QN(n1641) );
  NOR2X1 U2704 ( .IN1(reset), .IN2(n3176), .QN(n1642) );
  NOR2X1 U2705 ( .IN1(reset), .IN2(n3178), .QN(n1643) );
  NOR2X1 U2706 ( .IN1(reset), .IN2(n3144), .QN(n1618) );
  NOR2X1 U2707 ( .IN1(reset), .IN2(n3147), .QN(n1624) );
  NOR2X1 U2708 ( .IN1(reset), .IN2(n3149), .QN(n1625) );
  NOR2X1 U2709 ( .IN1(reset), .IN2(n3189), .QN(n1635) );
  NOR2X1 U2710 ( .IN1(reset), .IN2(n3153), .QN(n1620) );
  NOR2X1 U2711 ( .IN1(reset), .IN2(n3154), .QN(n1621) );
  NOR2X1 U2712 ( .IN1(reset), .IN2(n3155), .QN(n1626) );
  NOR2X1 U2713 ( .IN1(reset), .IN2(n3157), .QN(n1627) );
  NOR2X1 U2714 ( .IN1(reset), .IN2(n3146), .QN(n1619) );
  NOR2X1 U2715 ( .IN1(reset), .IN2(n3158), .QN(n1622) );
  NOR2X1 U2716 ( .IN1(reset), .IN2(n3159), .QN(n1628) );
  NOR2X1 U2717 ( .IN1(reset), .IN2(n3160), .QN(n1629) );
  NOR2X1 U2718 ( .IN1(reset), .IN2(n3161), .QN(n1637) );
  NOR2X1 U2719 ( .IN1(reset), .IN2(n3163), .QN(n1638) );
  NOR2X1 U2720 ( .IN1(reset), .IN2(n3181), .QN(n1634) );
  NOR2X1 U2721 ( .IN1(reset), .IN2(n3184), .QN(n1644) );
  NOR2X1 U2722 ( .IN1(reset), .IN2(n3187), .QN(n1645) );
  NOR2X1 U2723 ( .IN1(reset), .IN2(n3192), .QN(n1636) );
  IBUFFX4 U2724 ( .INP(search_data[24]), .ZN(n1726) );
  IBUFFX4 U2725 ( .INP(search_data[25]), .ZN(n1727) );
  NAND2X1 U2726 ( .IN1(n3123), .IN2(n3122), .QN(n3096) );
  NAND2X1 U2727 ( .IN1(n3114), .IN2(n3113), .QN(n3091) );
  NAND2X1 U2728 ( .IN1(n3088), .IN2(n3123), .QN(n2923) );
  NOR2X0 U2729 ( .IN1(n3188), .IN2(n3185), .QN(n3181) );
  NOR2X0 U2730 ( .IN1(n3188), .IN2(n3175), .QN(n3171) );
  NOR2X0 U2731 ( .IN1(n3177), .IN2(n3190), .QN(n3158) );
  NOR2X0 U2732 ( .IN1(n3188), .IN2(n3148), .QN(n3144) );
  NOR2X0 U2733 ( .IN1(n3183), .IN2(n3175), .QN(n3174) );
  NOR2X0 U2734 ( .IN1(n3186), .IN2(n3162), .QN(n3163) );
  NOR2X0 U2735 ( .IN1(n3190), .IN2(n3156), .QN(n3154) );
  NOR2X0 U2736 ( .IN1(n3183), .IN2(n3185), .QN(n3184) );
  NOR2X0 U2737 ( .IN1(n3191), .IN2(n3190), .QN(n3192) );
  NOR2X0 U2738 ( .IN1(n3186), .IN2(n3168), .QN(n3169) );
  NOR2X0 U2739 ( .IN1(n3183), .IN2(n3162), .QN(n3161) );
  NOR2X0 U2740 ( .IN1(n3148), .IN2(n3190), .QN(n3146) );
  NOR2X0 U2741 ( .IN1(n3186), .IN2(n3185), .QN(n3187) );
  NOR2X0 U2742 ( .IN1(n3186), .IN2(n3148), .QN(n3149) );
  NOR2X0 U2743 ( .IN1(n3186), .IN2(n3175), .QN(n3176) );
  NOR2X0 U2744 ( .IN1(n3191), .IN2(n3186), .QN(n3143) );
  NOR2X0 U2745 ( .IN1(n3190), .IN2(n3162), .QN(n3160) );
  NOR2X0 U2746 ( .IN1(n3188), .IN2(n3156), .QN(n3153) );
  NOR2X0 U2747 ( .IN1(n3177), .IN2(n3183), .QN(n3173) );
  NOR2X0 U2748 ( .IN1(n3190), .IN2(n3185), .QN(n3182) );
  NOR2X0 U2749 ( .IN1(n3183), .IN2(n3168), .QN(n3167) );
  NOR2X0 U2750 ( .IN1(n3188), .IN2(n3191), .QN(n3189) );
  NOR2X0 U2751 ( .IN1(n3177), .IN2(n3186), .QN(n3178) );
  NOR2X0 U2752 ( .IN1(n3188), .IN2(n3168), .QN(n3165) );
  NOR2X0 U2753 ( .IN1(n3183), .IN2(n3148), .QN(n3147) );
  NOR2X0 U2754 ( .IN1(n3190), .IN2(n3168), .QN(n3166) );
  NOR2X0 U2755 ( .IN1(n3186), .IN2(n3156), .QN(n3157) );
  NOR2X0 U2756 ( .IN1(n3188), .IN2(n3177), .QN(n3141) );
  NOR2X0 U2757 ( .IN1(n3183), .IN2(n3156), .QN(n3155) );
  NOR2X0 U2758 ( .IN1(n3188), .IN2(n3162), .QN(n3159) );
  NOR2X0 U2759 ( .IN1(n3190), .IN2(n3175), .QN(n3172) );
  NOR2X0 U2760 ( .IN1(n3191), .IN2(n3183), .QN(n3142) );
  NOR2X0 U2761 ( .IN1(write_index[4]), .IN2(n3150), .QN(n3180) );
  NOR2X0 U2762 ( .IN1(n3151), .IN2(n3150), .QN(n3170) );
  NAND2X0 U2763 ( .IN1(write), .IN2(n1742), .QN(n3150) );
  NOR2X0 U2764 ( .IN1(write_index[3]), .IN2(n3164), .QN(n3179) );
  INVX0 U2765 ( .INP(search), .ZN(n1611) );
  NOR2X0 U2766 ( .IN1(write_index[2]), .IN2(write_index[3]), .QN(n3152) );
  NOR4X0 U2767 ( .IN1(n2605), .IN2(n2604), .IN3(n1611), .IN4(n2603), .QN(n2629) );
  NAND2X1 U2768 ( .IN1(n3170), .IN2(n3179), .QN(n3162) );
  NAND2X1 U2769 ( .IN1(n3180), .IN2(n3179), .QN(n3185) );
  NAND2X1 U2770 ( .IN1(n3180), .IN2(n3152), .QN(n3177) );
  NAND2X1 U2771 ( .IN1(n3152), .IN2(n3170), .QN(n3156) );
  MUX21X1 U2772 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[25][24] ), .Q(n2734) );
  OR2X1 U2773 ( .IN1(n3145), .IN2(write_index[1]), .Q(n3190) );
  NAND2X1 U2774 ( .IN1(write_index[1]), .IN2(n3145), .QN(n3183) );
  INVX0 U2775 ( .INP(write_index[0]), .ZN(n3145) );
  INVX0 U2776 ( .INP(write_index[4]), .ZN(n3151) );
  NAND2X1 U2777 ( .IN1(write_index[1]), .IN2(write_index[0]), .QN(n3186) );
  INVX0 U2778 ( .INP(reset), .ZN(n1743) );
  OR2X1 U2779 ( .IN1(write_index[1]), .IN2(write_index[0]), .Q(n3188) );
  INVX0 U2780 ( .INP(write_index[2]), .ZN(n3164) );
  NAND2X0 U2781 ( .IN1(n1648), .IN2(n2840), .QN(n3012) );
  NAND2X0 U2782 ( .IN1(n3070), .IN2(n3069), .QN(n3107) );
  NOR2X0 U2783 ( .IN1(reset), .IN2(n3141), .QN(n1617) );
  NOR2X0 U2784 ( .IN1(reset), .IN2(n3182), .QN(n1616) );
  NOR2X0 U2785 ( .IN1(reset), .IN2(n3142), .QN(n1614) );
  NOR2X0 U2786 ( .IN1(reset), .IN2(n3173), .QN(n1615) );
  NOR4X0 U2787 ( .IN1(n2587), .IN2(n2586), .IN3(n2585), .IN4(n2584), .QN(n2590) );
  AND2X1 U2788 ( .IN1(n2589), .IN2(n2588), .Q(n1613) );
  NAND3X0 U2789 ( .IN1(write_index[2]), .IN2(write_index[3]), .IN3(n3170), 
        .QN(n3175) );
  NAND3X0 U2790 ( .IN1(n3180), .IN2(write_index[3]), .IN3(n3164), .QN(n3191)
         );
  NAND3X0 U2791 ( .IN1(n3180), .IN2(write_index[2]), .IN3(write_index[3]), 
        .QN(n3148) );
  NAND3X0 U2792 ( .IN1(write_index[3]), .IN2(n3170), .IN3(n3164), .QN(n3168)
         );
  AO221X1 U2793 ( .IN1(n1682), .IN2(\read_value_mux[31][7] ), .IN3(n1674), 
        .IN4(\read_value_mux[31][4] ), .IN5(n2594), .Q(n2632) );
  MUX21X1 U2794 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[31][25] ), .Q(n2599) );
  MUX21X1 U2795 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[29][23] ), .Q(n2575) );
  INVX0 U2796 ( .INP(reset), .ZN(n1742) );
  NAND2X0 U2797 ( .IN1(n3079), .IN2(n3078), .QN(n3109) );
  AND2X1 U2798 ( .IN1(n3076), .IN2(n3075), .Q(n1612) );
  IBUFFX32 U2799 ( .INP(search_data[23]), .ZN(n1725) );
  NAND2X0 U2800 ( .IN1(n3111), .IN2(n3110), .QN(n3081) );
  NAND3X1 U2801 ( .IN1(n3112), .IN2(n3111), .IN3(n3110), .QN(n3129) );
  IBUFFX4 U2802 ( .INP(search_data[28]), .ZN(n1733) );
  INVX0 U2803 ( .INP(search_data[26]), .ZN(n1728) );
  INVX0 U2804 ( .INP(search_data[16]), .ZN(n1708) );
  INVX0 U2805 ( .INP(search_data[13]), .ZN(n1700) );
  INVX0 U2806 ( .INP(search_data[19]), .ZN(n1716) );
  INVX0 U2807 ( .INP(search_data[15]), .ZN(n1705) );
  NAND2X1 U2808 ( .IN1(n3103), .IN2(n3102), .QN(n3137) );
  NAND2X1 U2809 ( .IN1(n3131), .IN2(n3130), .QN(n3134) );
  NAND2X1 U2810 ( .IN1(n3128), .IN2(n3127), .QN(n3135) );
  NAND2X1 U2811 ( .IN1(n3095), .IN2(n3094), .QN(n3106) );
  NAND2X1 U2812 ( .IN1(n3067), .IN2(n3066), .QN(n3108) );
  MUX21X1 U2813 ( .IN1(n1700), .IN2(search_data[13]), .S(
        \read_value_mux[0][13] ), .Q(n1786) );
  MUX21X1 U2814 ( .IN1(n1692), .IN2(search_data[10]), .S(
        \read_value_mux[25][10] ), .Q(n2743) );
  MUX21X1 U2815 ( .IN1(n1673), .IN2(search_data[4]), .S(
        \read_value_mux[29][4] ), .Q(n2582) );
  MUX21X1 U2816 ( .IN1(n1688), .IN2(search_data[9]), .S(
        \read_value_mux[29][9] ), .Q(n2577) );
  MUX21X1 U2817 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[29][24] ), .Q(n2568) );
  MUX21X1 U2818 ( .IN1(n1698), .IN2(search_data[13]), .S(
        \read_value_mux[28][13] ), .Q(n2685) );
  INVX0 U2819 ( .INP(search_data[7]), .ZN(n1683) );
  MUX21X1 U2820 ( .IN1(n1694), .IN2(search_data[11]), .S(
        \read_value_mux[31][11] ), .Q(n2620) );
  MUX21X1 U2821 ( .IN1(n1684), .IN2(search_data[8]), .S(
        \read_value_mux[31][8] ), .Q(n2615) );
  MUX21X1 U2822 ( .IN1(n1692), .IN2(search_data[10]), .S(
        \read_value_mux[31][10] ), .Q(n2611) );
  MUX21X1 U2823 ( .IN1(n1729), .IN2(search_data[26]), .S(
        \read_value_mux[31][26] ), .Q(n2608) );
  MUX21X1 U2824 ( .IN1(n1699), .IN2(search_data[13]), .S(
        \read_value_mux[30][13] ), .Q(n2662) );
  INVX0 U2825 ( .INP(search_data[5]), .ZN(n1675) );
  INVX0 U2826 ( .INP(search_data[14]), .ZN(n1702) );
  INVX0 U2827 ( .INP(search_data[26]), .ZN(n1729) );
  INVX0 U2828 ( .INP(search_data[8]), .ZN(n1684) );
  INVX0 U2829 ( .INP(search_data[12]), .ZN(n1697) );
  INVX0 U2830 ( .INP(search_data[30]), .ZN(n1737) );
  INVX0 U2831 ( .INP(search_data[3]), .ZN(n1669) );
  INVX0 U2832 ( .INP(search_data[6]), .ZN(n1678) );
  INVX0 U2833 ( .INP(search_data[29]), .ZN(n1734) );
  INVX0 U2834 ( .INP(search_data[13]), .ZN(n1698) );
  INVX0 U2835 ( .INP(search_data[21]), .ZN(n1719) );
  INVX0 U2836 ( .INP(search_data[9]), .ZN(n1687) );
  INVX0 U2837 ( .INP(search_data[22]), .ZN(n1722) );
  INVX0 U2838 ( .INP(search_data[5]), .ZN(n1677) );
  INVX0 U2839 ( .INP(search_data[2]), .ZN(n1666) );
  INVX0 U2840 ( .INP(search_data[16]), .ZN(n1707) );
  INVX0 U2841 ( .INP(search_data[13]), .ZN(n1699) );
  INVX0 U2842 ( .INP(search_data[1]), .ZN(n1664) );
  INVX0 U2843 ( .INP(search_data[18]), .ZN(n1713) );
  INVX0 U2844 ( .INP(search_data[17]), .ZN(n1710) );
  INVX0 U2845 ( .INP(search_data[6]), .ZN(n1679) );
  INVX0 U2846 ( .INP(search_data[9]), .ZN(n1688) );
  INVX0 U2847 ( .INP(search_data[4]), .ZN(n1673) );
  INVX0 U2848 ( .INP(search_data[22]), .ZN(n1723) );
  INVX0 U2849 ( .INP(search_data[14]), .ZN(n1701) );
  INVX0 U2850 ( .INP(search_data[0]), .ZN(n1661) );
  MUX21X1 U2851 ( .IN1(n1700), .IN2(search_data[13]), .S(
        \read_value_mux[7][13] ), .Q(n1942) );
  INVX0 U2852 ( .INP(search_data[19]), .ZN(n1717) );
  INVX0 U2853 ( .INP(search_data[11]), .ZN(n1694) );
  INVX0 U2854 ( .INP(search_data[29]), .ZN(n1735) );
  INVX0 U2855 ( .INP(search_data[0]), .ZN(n1662) );
  MUX21X1 U2856 ( .IN1(n1700), .IN2(search_data[13]), .S(
        \read_value_mux[6][13] ), .Q(n1976) );
  INVX0 U2857 ( .INP(search_data[18]), .ZN(n1712) );
  INVX0 U2858 ( .INP(search_data[15]), .ZN(n1706) );
  INVX0 U2859 ( .INP(search_data[10]), .ZN(n1692) );
  INVX0 U2860 ( .INP(search_data[21]), .ZN(n1721) );
  INVX0 U2861 ( .INP(search_data[2]), .ZN(n1667) );
  INVX0 U2862 ( .INP(search_data[8]), .ZN(n1686) );
  INVX0 U2863 ( .INP(search_data[27]), .ZN(n1732) );
  INVX0 U2864 ( .INP(search_data[17]), .ZN(n1709) );
  INVX0 U2865 ( .INP(search_data[4]), .ZN(n1672) );
  INVX0 U2866 ( .INP(search_data[31]), .ZN(n1741) );
  INVX0 U2867 ( .INP(search_data[11]), .ZN(n1695) );
  MUX21X1 U2868 ( .IN1(n1700), .IN2(search_data[13]), .S(
        \read_value_mux[5][13] ), .Q(n1890) );
  INVX0 U2869 ( .INP(search_data[30]), .ZN(n1739) );
  INVX0 U2870 ( .INP(search_data[27]), .ZN(n1731) );
  INVX0 U2871 ( .INP(search_data[7]), .ZN(n1682) );
  INVX0 U2872 ( .INP(search_data[19]), .ZN(n1715) );
  INVX0 U2873 ( .INP(search_data[1]), .ZN(n1663) );
  INVX0 U2874 ( .INP(search_data[27]), .ZN(n1730) );
  NBUFFX2 U2875 ( .INP(search_data[10]), .Z(n1690) );
  INVX0 U2876 ( .INP(search_data[1]), .ZN(n1665) );
  INVX0 U2877 ( .INP(search_data[21]), .ZN(n1720) );
  INVX0 U2878 ( .INP(search_data[8]), .ZN(n1685) );
  NBUFFX2 U2879 ( .INP(search_data[15]), .Z(n1704) );
  INVX0 U2880 ( .INP(search_data[18]), .ZN(n1714) );
  INVX0 U2881 ( .INP(search_data[0]), .ZN(n1660) );
  INVX0 U2882 ( .INP(search_data[30]), .ZN(n1738) );
  INVX0 U2883 ( .INP(search_data[17]), .ZN(n1711) );
  MUX21X1 U2884 ( .IN1(n1700), .IN2(search_data[13]), .S(
        \read_value_mux[4][13] ), .Q(n2000) );
  INVX0 U2885 ( .INP(search_data[5]), .ZN(n1676) );
  INVX0 U2886 ( .INP(search_data[3]), .ZN(n1670) );
  INVX0 U2887 ( .INP(search), .ZN(n1659) );
  INVX0 U2888 ( .INP(search_data[31]), .ZN(n1740) );
  INVX0 U2889 ( .INP(search_data[22]), .ZN(n1724) );
  INVX0 U2890 ( .INP(search_data[2]), .ZN(n1668) );
  INVX0 U2891 ( .INP(search_data[4]), .ZN(n1674) );
  INVX0 U2892 ( .INP(search_data[12]), .ZN(n1696) );
  INVX0 U2893 ( .INP(search_data[9]), .ZN(n1689) );
  INVX0 U2894 ( .INP(search_data[14]), .ZN(n1703) );
  INVX0 U2895 ( .INP(search_data[29]), .ZN(n1736) );
  INVX0 U2896 ( .INP(search_data[11]), .ZN(n1693) );
  INVX0 U2897 ( .INP(search_data[7]), .ZN(n1681) );
  INVX0 U2898 ( .INP(search_data[6]), .ZN(n1680) );
  OR3X1 U2899 ( .IN1(n2631), .IN2(n2632), .IN3(n2633), .Q(n1646) );
  OR2X1 U2900 ( .IN1(n3118), .IN2(n3120), .Q(n1647) );
  AND2X1 U2901 ( .IN1(n3082), .IN2(n3008), .Q(n1648) );
  NAND3X0 U2902 ( .IN1(n3094), .IN2(n3012), .IN3(n3011), .QN(n1654) );
  AND4X1 U2903 ( .IN1(n3055), .IN2(n3095), .IN3(n3060), .IN4(n3057), .Q(n1655)
         );
  NOR2X0 U2904 ( .IN1(n3101), .IN2(n1647), .QN(search_index[1]) );
  OAI221X1 U2905 ( .IN1(search_data[3]), .IN2(n1656), .IN3(n1657), .IN4(
        search_data[23]), .IN5(n1658), .QN(n2633) );
  OA22X1 U2906 ( .IN1(n1671), .IN2(\read_value_mux[31][3] ), .IN3(n1725), 
        .IN4(\read_value_mux[31][23] ), .Q(n1658) );
  INVX0 U2907 ( .INP(search_data[3]), .ZN(n1671) );
  OR2X1 U2908 ( .IN1(n2630), .IN2(n1646), .Q(n3075) );
  MUX41X1 U2909 ( .IN1(\words[0]/valid_o ), .IN3(\words[1]/valid_o ), .IN2(
        \words[2]/valid_o ), .IN4(\words[3]/valid_o ), .S0(read_index[0]), 
        .S1(read_index[1]), .Q(n1747) );
  MUX41X1 U2910 ( .IN1(\words[8]/valid_o ), .IN3(\words[9]/valid_o ), .IN2(
        \words[10]/valid_o ), .IN4(\words[11]/valid_o ), .S0(read_index[0]), 
        .S1(read_index[1]), .Q(n1746) );
  MUX41X1 U2911 ( .IN1(\words[4]/valid_o ), .IN3(\words[5]/valid_o ), .IN2(
        \words[6]/valid_o ), .IN4(\words[7]/valid_o ), .S0(read_index[0]), 
        .S1(read_index[1]), .Q(n1745) );
  MUX41X1 U2912 ( .IN1(\words[12]/valid_o ), .IN3(\words[13]/valid_o ), .IN2(
        \words[14]/valid_o ), .IN4(\words[15]/valid_o ), .S0(read_index[0]), 
        .S1(read_index[1]), .Q(n1744) );
  MUX41X1 U2913 ( .IN1(n1747), .IN3(n1746), .IN2(n1745), .IN4(n1744), .S0(
        read_index[3]), .S1(read_index[2]), .Q(n1754) );
  INVX0 U2914 ( .INP(read_index[4]), .ZN(n1753) );
  MUX41X1 U2915 ( .IN1(\words[16]/valid_o ), .IN3(\words[17]/valid_o ), .IN2(
        \words[18]/valid_o ), .IN4(\words[19]/valid_o ), .S0(read_index[0]), 
        .S1(read_index[1]), .Q(n1751) );
  MUX41X1 U2916 ( .IN1(\words[24]/valid_o ), .IN3(\words[25]/valid_o ), .IN2(
        \words[26]/valid_o ), .IN4(\words[27]/valid_o ), .S0(read_index[0]), 
        .S1(read_index[1]), .Q(n1750) );
  MUX41X1 U2917 ( .IN1(\words[20]/valid_o ), .IN3(\words[21]/valid_o ), .IN2(
        \words[22]/valid_o ), .IN4(\words[23]/valid_o ), .S0(read_index[0]), 
        .S1(read_index[1]), .Q(n1749) );
  MUX41X1 U2918 ( .IN1(\words[28]/valid_o ), .IN3(\words[29]/valid_o ), .IN2(
        \words[30]/valid_o ), .IN4(\words[31]/valid_o ), .S0(read_index[0]), 
        .S1(read_index[1]), .Q(n1748) );
  MUX41X1 U2919 ( .IN1(n1751), .IN3(n1750), .IN2(n1749), .IN4(n1748), .S0(
        read_index[3]), .S1(read_index[2]), .Q(n1752) );
  OA221X1 U2920 ( .IN1(read_index[4]), .IN2(n1754), .IN3(n1753), .IN4(n1752), 
        .IN5(read), .Q(read_valid) );
  MUX21X1 U2921 ( .IN1(search_data[26]), .IN2(n1728), .S(
        \read_value_mux[0][26] ), .Q(n1763) );
  MUX21X1 U2922 ( .IN1(search_data[7]), .IN2(n1681), .S(\read_value_mux[0][7] ), .Q(n1762) );
  OAI22X1 U2923 ( .IN1(\read_value_mux[0][6] ), .IN2(n1680), .IN3(n1713), 
        .IN4(\read_value_mux[0][18] ), .QN(n1755) );
  AO221X1 U2924 ( .IN1(n1680), .IN2(\read_value_mux[0][6] ), .IN3(n1712), 
        .IN4(\read_value_mux[0][18] ), .IN5(n1755), .Q(n1761) );
  MUX21X1 U2925 ( .IN1(n1716), .IN2(search_data[19]), .S(
        \read_value_mux[0][19] ), .Q(n1759) );
  MUX21X1 U2926 ( .IN1(n1666), .IN2(search_data[2]), .S(\read_value_mux[0][2] ), .Q(n1757) );
  MUX21X1 U2927 ( .IN1(n1709), .IN2(search_data[17]), .S(
        \read_value_mux[0][17] ), .Q(n1756) );
  NAND4X0 U2928 ( .IN1(n1759), .IN2(n1758), .IN3(n1757), .IN4(n1756), .QN(
        n1760) );
  NOR4X0 U2929 ( .IN1(n1763), .IN2(n1762), .IN3(n1761), .IN4(n1760), .QN(n1795) );
  MUX21X1 U2930 ( .IN1(n1669), .IN2(search_data[3]), .S(\read_value_mux[0][3] ), .Q(n1764) );
  OA221X1 U2931 ( .IN1(search_data[27]), .IN2(n1650), .IN3(n1732), .IN4(
        \read_value_mux[0][27] ), .IN5(n1764), .Q(n1794) );
  MUX21X1 U2932 ( .IN1(search_data[15]), .IN2(n1705), .S(
        \read_value_mux[0][15] ), .Q(n1771) );
  MUX21X1 U2933 ( .IN1(search_data[9]), .IN2(n1687), .S(\read_value_mux[0][9] ), .Q(n1770) );
  MUX21X1 U2934 ( .IN1(n1693), .IN2(search_data[11]), .S(
        \read_value_mux[0][11] ), .Q(n1768) );
  MUX21X1 U2935 ( .IN1(n1672), .IN2(search_data[4]), .S(\read_value_mux[0][4] ), .Q(n1767) );
  MUX21X1 U2936 ( .IN1(n1737), .IN2(search_data[30]), .S(
        \read_value_mux[0][30] ), .Q(n1766) );
  MUX21X1 U2937 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[0][25] ), .Q(n1765) );
  NAND4X0 U2938 ( .IN1(n1768), .IN2(n1767), .IN3(n1766), .IN4(n1765), .QN(
        n1769) );
  NOR4X0 U2939 ( .IN1(n1771), .IN2(n1770), .IN3(n1659), .IN4(n1769), .QN(n1793) );
  MUX21X1 U2940 ( .IN1(n1734), .IN2(search_data[29]), .S(
        \read_value_mux[0][29] ), .Q(n1775) );
  MUX21X1 U2941 ( .IN1(n1691), .IN2(n1690), .S(\read_value_mux[0][10] ), .Q(
        n1774) );
  MUX21X1 U2942 ( .IN1(n1718), .IN2(search_data[20]), .S(
        \read_value_mux[0][20] ), .Q(n1773) );
  MUX21X1 U2943 ( .IN1(n1684), .IN2(search_data[8]), .S(\read_value_mux[0][8] ), .Q(n1772) );
  NAND4X0 U2944 ( .IN1(n1775), .IN2(n1774), .IN3(n1773), .IN4(n1772), .QN(
        n1791) );
  MUX21X1 U2945 ( .IN1(n1701), .IN2(search_data[14]), .S(
        \read_value_mux[0][14] ), .Q(n1779) );
  MUX21X1 U2946 ( .IN1(n1660), .IN2(search_data[0]), .S(\read_value_mux[0][0] ), .Q(n1778) );
  MUX21X1 U2947 ( .IN1(n1675), .IN2(search_data[5]), .S(\read_value_mux[0][5] ), .Q(n1777) );
  MUX21X1 U2948 ( .IN1(n1708), .IN2(search_data[16]), .S(
        \read_value_mux[0][16] ), .Q(n1776) );
  NAND4X0 U2949 ( .IN1(n1779), .IN2(n1778), .IN3(n1777), .IN4(n1776), .QN(
        n1790) );
  MUX21X1 U2950 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[0][23] ), .Q(n1783) );
  MUX21X1 U2951 ( .IN1(n1740), .IN2(search_data[31]), .S(
        \read_value_mux[0][31] ), .Q(n1782) );
  MUX21X1 U2952 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[0][24] ), .Q(n1781) );
  MUX21X1 U2953 ( .IN1(n1665), .IN2(search_data[1]), .S(\read_value_mux[0][1] ), .Q(n1780) );
  NAND4X0 U2954 ( .IN1(n1783), .IN2(n1782), .IN3(n1781), .IN4(n1780), .QN(
        n1789) );
  MUX21X1 U2955 ( .IN1(n1697), .IN2(search_data[12]), .S(
        \read_value_mux[0][12] ), .Q(n1787) );
  MUX21X1 U2956 ( .IN1(n1719), .IN2(search_data[21]), .S(
        \read_value_mux[0][21] ), .Q(n1785) );
  MUX21X1 U2957 ( .IN1(n1722), .IN2(search_data[22]), .S(
        \read_value_mux[0][22] ), .Q(n1784) );
  NAND4X0 U2958 ( .IN1(n1787), .IN2(n1786), .IN3(n1785), .IN4(n1784), .QN(
        n1788) );
  NOR4X0 U2959 ( .IN1(n1791), .IN2(n1790), .IN3(n1789), .IN4(n1788), .QN(n1792) );
  NAND4X0 U2960 ( .IN1(n1795), .IN2(n1794), .IN3(n1793), .IN4(n1792), .QN(
        n3056) );
  MUX21X1 U2961 ( .IN1(search_data[12]), .IN2(n1696), .S(
        \read_value_mux[2][12] ), .Q(n1804) );
  MUX21X1 U2962 ( .IN1(search_data[0]), .IN2(n1662), .S(\read_value_mux[2][0] ), .Q(n1803) );
  OAI22X1 U2963 ( .IN1(\read_value_mux[2][13] ), .IN2(n1700), .IN3(n1706), 
        .IN4(\read_value_mux[2][15] ), .QN(n1796) );
  AO221X1 U2964 ( .IN1(n1700), .IN2(\read_value_mux[2][13] ), .IN3(n1706), 
        .IN4(\read_value_mux[2][15] ), .IN5(n1796), .Q(n1802) );
  MUX21X1 U2965 ( .IN1(n1687), .IN2(search_data[9]), .S(\read_value_mux[2][9] ), .Q(n1800) );
  MUX21X1 U2966 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[2][25] ), .Q(n1799) );
  MUX21X1 U2967 ( .IN1(n1667), .IN2(search_data[2]), .S(\read_value_mux[2][2] ), .Q(n1798) );
  MUX21X1 U2968 ( .IN1(n1710), .IN2(search_data[17]), .S(
        \read_value_mux[2][17] ), .Q(n1797) );
  NAND4X0 U2969 ( .IN1(n1800), .IN2(n1799), .IN3(n1798), .IN4(n1797), .QN(
        n1801) );
  NOR4X0 U2970 ( .IN1(n1804), .IN2(n1803), .IN3(n1802), .IN4(n1801), .QN(n1836) );
  MUX21X1 U2971 ( .IN1(n1739), .IN2(search_data[30]), .S(
        \read_value_mux[2][30] ), .Q(n1805) );
  OA221X1 U2972 ( .IN1(search_data[5]), .IN2(n1651), .IN3(n1677), .IN4(
        \read_value_mux[2][5] ), .IN5(n1805), .Q(n1835) );
  MUX21X1 U2973 ( .IN1(search_data[27]), .IN2(n1730), .S(
        \read_value_mux[2][27] ), .Q(n1812) );
  MUX21X1 U2974 ( .IN1(search_data[19]), .IN2(n1717), .S(
        \read_value_mux[2][19] ), .Q(n1811) );
  MUX21X1 U2975 ( .IN1(n1685), .IN2(search_data[8]), .S(\read_value_mux[2][8] ), .Q(n1809) );
  MUX21X1 U2976 ( .IN1(n1724), .IN2(search_data[22]), .S(
        \read_value_mux[2][22] ), .Q(n1808) );
  MUX21X1 U2977 ( .IN1(n1673), .IN2(search_data[4]), .S(\read_value_mux[2][4] ), .Q(n1807) );
  MUX21X1 U2978 ( .IN1(n1681), .IN2(search_data[7]), .S(\read_value_mux[2][7] ), .Q(n1806) );
  NAND4X0 U2979 ( .IN1(n1809), .IN2(n1808), .IN3(n1807), .IN4(n1806), .QN(
        n1810) );
  NOR4X0 U2980 ( .IN1(n1812), .IN2(n1811), .IN3(n1659), .IN4(n1810), .QN(n1834) );
  MUX21X1 U2981 ( .IN1(n1721), .IN2(search_data[21]), .S(
        \read_value_mux[2][21] ), .Q(n1816) );
  MUX21X1 U2982 ( .IN1(n1718), .IN2(search_data[20]), .S(
        \read_value_mux[2][20] ), .Q(n1815) );
  MUX21X1 U2983 ( .IN1(n1735), .IN2(search_data[29]), .S(
        \read_value_mux[2][29] ), .Q(n1813) );
  NAND4X0 U2984 ( .IN1(n1816), .IN2(n1815), .IN3(n1814), .IN4(n1813), .QN(
        n1832) );
  MUX21X1 U2985 ( .IN1(n1702), .IN2(search_data[14]), .S(
        \read_value_mux[2][14] ), .Q(n1820) );
  MUX21X1 U2986 ( .IN1(n1680), .IN2(search_data[6]), .S(\read_value_mux[2][6] ), .Q(n1819) );
  MUX21X1 U2987 ( .IN1(n1670), .IN2(search_data[3]), .S(\read_value_mux[2][3] ), .Q(n1818) );
  MUX21X1 U2988 ( .IN1(n1707), .IN2(search_data[16]), .S(
        \read_value_mux[2][16] ), .Q(n1817) );
  NAND4X0 U2989 ( .IN1(n1820), .IN2(n1819), .IN3(n1818), .IN4(n1817), .QN(
        n1831) );
  MUX21X1 U2990 ( .IN1(n1714), .IN2(search_data[18]), .S(
        \read_value_mux[2][18] ), .Q(n1824) );
  MUX21X1 U2991 ( .IN1(n1740), .IN2(search_data[31]), .S(
        \read_value_mux[2][31] ), .Q(n1823) );
  MUX21X1 U2992 ( .IN1(n1695), .IN2(search_data[11]), .S(
        \read_value_mux[2][11] ), .Q(n1822) );
  MUX21X1 U2993 ( .IN1(n1665), .IN2(search_data[1]), .S(\read_value_mux[2][1] ), .Q(n1821) );
  NAND4X0 U2994 ( .IN1(n1824), .IN2(n1823), .IN3(n1822), .IN4(n1821), .QN(
        n1830) );
  MUX21X1 U2995 ( .IN1(n1728), .IN2(search_data[26]), .S(
        \read_value_mux[2][26] ), .Q(n1828) );
  MUX21X1 U2996 ( .IN1(n1692), .IN2(n1690), .S(\read_value_mux[2][10] ), .Q(
        n1827) );
  MUX21X1 U2997 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[2][23] ), .Q(n1826) );
  MUX21X1 U2998 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[2][24] ), .Q(n1825) );
  NAND4X0 U2999 ( .IN1(n1828), .IN2(n1827), .IN3(n1826), .IN4(n1825), .QN(
        n1829) );
  NOR4X0 U3000 ( .IN1(n1832), .IN2(n1831), .IN3(n1830), .IN4(n1829), .QN(n1833) );
  NAND4X0 U3001 ( .IN1(n1836), .IN2(n1835), .IN3(n1834), .IN4(n1833), .QN(
        n3013) );
  OAI22X1 U3002 ( .IN1(\read_value_mux[3][15] ), .IN2(n1706), .IN3(n1714), 
        .IN4(\read_value_mux[3][18] ), .QN(n1837) );
  AO221X1 U3003 ( .IN1(n1706), .IN2(\read_value_mux[3][15] ), .IN3(n1713), 
        .IN4(\read_value_mux[3][18] ), .IN5(n1837), .Q(n1870) );
  OAI22X1 U3004 ( .IN1(\read_value_mux[3][0] ), .IN2(n1660), .IN3(n1689), 
        .IN4(\read_value_mux[3][9] ), .QN(n1838) );
  AO221X1 U3005 ( .IN1(n1661), .IN2(\read_value_mux[3][0] ), .IN3(n1689), 
        .IN4(\read_value_mux[3][9] ), .IN5(n1838), .Q(n1869) );
  MUX21X1 U3006 ( .IN1(n1711), .IN2(search_data[17]), .S(
        \read_value_mux[3][17] ), .Q(n1842) );
  MUX21X1 U3007 ( .IN1(n1665), .IN2(search_data[1]), .S(\read_value_mux[3][1] ), .Q(n1841) );
  MUX21X1 U3008 ( .IN1(n1730), .IN2(search_data[27]), .S(
        \read_value_mux[3][27] ), .Q(n1840) );
  MUX21X1 U3009 ( .IN1(n1721), .IN2(search_data[21]), .S(
        \read_value_mux[3][21] ), .Q(n1839) );
  NAND4X0 U3010 ( .IN1(n1842), .IN2(n1841), .IN3(n1840), .IN4(n1839), .QN(
        n1868) );
  MUX21X1 U3011 ( .IN1(n1695), .IN2(search_data[11]), .S(
        \read_value_mux[3][11] ), .Q(n1846) );
  MUX21X1 U3012 ( .IN1(n1691), .IN2(n1690), .S(\read_value_mux[3][10] ), .Q(
        n1845) );
  MUX21X1 U3013 ( .IN1(n1718), .IN2(search_data[20]), .S(
        \read_value_mux[3][20] ), .Q(n1844) );
  MUX21X1 U3014 ( .IN1(n1739), .IN2(search_data[30]), .S(
        \read_value_mux[3][30] ), .Q(n1843) );
  NAND4X0 U3015 ( .IN1(n1846), .IN2(n1845), .IN3(n1844), .IN4(n1843), .QN(
        n1862) );
  MUX21X1 U3016 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[3][25] ), .Q(n1850) );
  MUX21X1 U3017 ( .IN1(n1671), .IN2(search_data[3]), .S(\read_value_mux[3][3] ), .Q(n1849) );
  MUX21X1 U3018 ( .IN1(n1680), .IN2(search_data[6]), .S(\read_value_mux[3][6] ), .Q(n1848) );
  MUX21X1 U3019 ( .IN1(n1696), .IN2(search_data[12]), .S(
        \read_value_mux[3][12] ), .Q(n1847) );
  NAND4X0 U3020 ( .IN1(n1850), .IN2(n1849), .IN3(n1848), .IN4(n1847), .QN(
        n1861) );
  MUX21X1 U3021 ( .IN1(n1728), .IN2(search_data[26]), .S(
        \read_value_mux[3][26] ), .Q(n1854) );
  MUX21X1 U3022 ( .IN1(n1708), .IN2(search_data[16]), .S(
        \read_value_mux[3][16] ), .Q(n1853) );
  MUX21X1 U3023 ( .IN1(n1724), .IN2(search_data[22]), .S(
        \read_value_mux[3][22] ), .Q(n1852) );
  MUX21X1 U3024 ( .IN1(n1668), .IN2(search_data[2]), .S(\read_value_mux[3][2] ), .Q(n1851) );
  NAND4X0 U3025 ( .IN1(n1854), .IN2(n1853), .IN3(n1852), .IN4(n1851), .QN(
        n1860) );
  MUX21X1 U3026 ( .IN1(n1686), .IN2(search_data[8]), .S(\read_value_mux[3][8] ), .Q(n1858) );
  MUX21X1 U3027 ( .IN1(n1674), .IN2(search_data[4]), .S(\read_value_mux[3][4] ), .Q(n1857) );
  MUX21X1 U3028 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[3][23] ), .Q(n1856) );
  MUX21X1 U3029 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[3][24] ), .Q(n1855) );
  NAND4X0 U3030 ( .IN1(n1858), .IN2(n1857), .IN3(n1856), .IN4(n1855), .QN(
        n1859) );
  NOR4X0 U3031 ( .IN1(n1862), .IN2(n1861), .IN3(n1860), .IN4(n1859), .QN(n1865) );
  MUX21X1 U3032 ( .IN1(n1682), .IN2(search_data[7]), .S(\read_value_mux[3][7] ), .Q(n1864) );
  MUX21X1 U3033 ( .IN1(n1736), .IN2(search_data[29]), .S(
        \read_value_mux[3][29] ), .Q(n1863) );
  NAND4X0 U3034 ( .IN1(n1866), .IN2(n1865), .IN3(n1864), .IN4(n1863), .QN(
        n1867) );
  NOR4X0 U3035 ( .IN1(n1870), .IN2(n1869), .IN3(n1868), .IN4(n1867), .QN(n3117) );
  MUX21X1 U3036 ( .IN1(search_data[1]), .IN2(n1663), .S(\read_value_mux[5][1] ), .Q(n1911) );
  MUX21X1 U3037 ( .IN1(search_data[19]), .IN2(n1715), .S(
        \read_value_mux[5][19] ), .Q(n1910) );
  AOI22X1 U3038 ( .IN1(n1733), .IN2(\read_value_mux[5][28] ), .IN3(n1708), 
        .IN4(\read_value_mux[5][16] ), .QN(n1871) );
  OA221X1 U3039 ( .IN1(n1733), .IN2(\read_value_mux[5][28] ), .IN3(n1708), 
        .IN4(\read_value_mux[5][16] ), .IN5(n1871), .Q(n1876) );
  AOI22X1 U3040 ( .IN1(n1724), .IN2(\read_value_mux[5][22] ), .IN3(n1726), 
        .IN4(\read_value_mux[5][24] ), .QN(n1872) );
  OA221X1 U3041 ( .IN1(n1724), .IN2(\read_value_mux[5][22] ), .IN3(n1726), 
        .IN4(\read_value_mux[5][24] ), .IN5(n1872), .Q(n1875) );
  MUX21X1 U3042 ( .IN1(n1728), .IN2(search_data[26]), .S(
        \read_value_mux[5][26] ), .Q(n1874) );
  MUX21X1 U3043 ( .IN1(n1705), .IN2(n1704), .S(\read_value_mux[5][15] ), .Q(
        n1873) );
  NAND4X0 U3044 ( .IN1(n1876), .IN2(n1875), .IN3(n1874), .IN4(n1873), .QN(
        n1909) );
  MUX21X1 U3045 ( .IN1(search_data[23]), .IN2(n1725), .S(
        \read_value_mux[5][23] ), .Q(n1883) );
  MUX21X1 U3046 ( .IN1(search_data[20]), .IN2(n1718), .S(
        \read_value_mux[5][20] ), .Q(n1882) );
  MUX21X1 U3047 ( .IN1(n1720), .IN2(search_data[21]), .S(
        \read_value_mux[5][21] ), .Q(n1880) );
  MUX21X1 U3048 ( .IN1(n1682), .IN2(search_data[7]), .S(\read_value_mux[5][7] ), .Q(n1879) );
  MUX21X1 U3049 ( .IN1(n1731), .IN2(search_data[27]), .S(
        \read_value_mux[5][27] ), .Q(n1878) );
  MUX21X1 U3050 ( .IN1(n1676), .IN2(search_data[5]), .S(\read_value_mux[5][5] ), .Q(n1877) );
  NAND4X0 U3051 ( .IN1(n1880), .IN2(n1879), .IN3(n1878), .IN4(n1877), .QN(
        n1881) );
  NOR4X0 U3052 ( .IN1(n1883), .IN2(n1882), .IN3(n1659), .IN4(n1881), .QN(n1907) );
  MUX21X1 U3053 ( .IN1(n1739), .IN2(search_data[30]), .S(
        \read_value_mux[5][30] ), .Q(n1887) );
  MUX21X1 U3054 ( .IN1(n1671), .IN2(search_data[3]), .S(\read_value_mux[5][3] ), .Q(n1886) );
  MUX21X1 U3055 ( .IN1(n1685), .IN2(search_data[8]), .S(\read_value_mux[5][8] ), .Q(n1885) );
  MUX21X1 U3056 ( .IN1(n1711), .IN2(search_data[17]), .S(
        \read_value_mux[5][17] ), .Q(n1884) );
  NAND4X0 U3057 ( .IN1(n1887), .IN2(n1886), .IN3(n1885), .IN4(n1884), .QN(
        n1903) );
  MUX21X1 U3058 ( .IN1(n1703), .IN2(search_data[14]), .S(
        \read_value_mux[5][14] ), .Q(n1891) );
  MUX21X1 U3059 ( .IN1(n1714), .IN2(search_data[18]), .S(
        \read_value_mux[5][18] ), .Q(n1889) );
  MUX21X1 U3060 ( .IN1(n1736), .IN2(search_data[29]), .S(
        \read_value_mux[5][29] ), .Q(n1888) );
  NAND4X0 U3061 ( .IN1(n1891), .IN2(n1890), .IN3(n1889), .IN4(n1888), .QN(
        n1902) );
  MUX21X1 U3062 ( .IN1(n1696), .IN2(search_data[12]), .S(
        \read_value_mux[5][12] ), .Q(n1895) );
  MUX21X1 U3063 ( .IN1(n1660), .IN2(search_data[0]), .S(\read_value_mux[5][0] ), .Q(n1894) );
  MUX21X1 U3064 ( .IN1(n1680), .IN2(search_data[6]), .S(\read_value_mux[5][6] ), .Q(n1893) );
  MUX21X1 U3065 ( .IN1(n1691), .IN2(n1690), .S(\read_value_mux[5][10] ), .Q(
        n1892) );
  NAND4X0 U3066 ( .IN1(n1895), .IN2(n1894), .IN3(n1893), .IN4(n1892), .QN(
        n1901) );
  MUX21X1 U3067 ( .IN1(n1668), .IN2(search_data[2]), .S(\read_value_mux[5][2] ), .Q(n1899) );
  MUX21X1 U3068 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[5][25] ), .Q(n1898) );
  MUX21X1 U3069 ( .IN1(n1695), .IN2(search_data[11]), .S(
        \read_value_mux[5][11] ), .Q(n1897) );
  MUX21X1 U3070 ( .IN1(n1674), .IN2(search_data[4]), .S(\read_value_mux[5][4] ), .Q(n1896) );
  NAND4X0 U3071 ( .IN1(n1899), .IN2(n1898), .IN3(n1897), .IN4(n1896), .QN(
        n1900) );
  NOR4X0 U3072 ( .IN1(n1903), .IN2(n1902), .IN3(n1901), .IN4(n1900), .QN(n1906) );
  MUX21X1 U3073 ( .IN1(n1689), .IN2(search_data[9]), .S(\read_value_mux[5][9] ), .Q(n1905) );
  MUX21X1 U3074 ( .IN1(n1741), .IN2(search_data[31]), .S(
        \read_value_mux[5][31] ), .Q(n1904) );
  NAND4X0 U3075 ( .IN1(n1907), .IN2(n1906), .IN3(n1905), .IN4(n1904), .QN(
        n1908) );
  NOR4X0 U3076 ( .IN1(n1911), .IN2(n1910), .IN3(n1909), .IN4(n1908), .QN(n3058) );
  MUX21X1 U3077 ( .IN1(search_data[26]), .IN2(n1728), .S(
        \read_value_mux[7][26] ), .Q(n1948) );
  MUX21X1 U3078 ( .IN1(n1690), .IN2(n1691), .S(\read_value_mux[7][10] ), .Q(
        n1947) );
  AOI22X1 U3079 ( .IN1(n1706), .IN2(\read_value_mux[7][15] ), .IN3(n1739), 
        .IN4(\read_value_mux[7][30] ), .QN(n1912) );
  OA221X1 U3080 ( .IN1(n1706), .IN2(\read_value_mux[7][15] ), .IN3(n1739), 
        .IN4(\read_value_mux[7][30] ), .IN5(n1912), .Q(n1917) );
  AOI22X1 U3081 ( .IN1(n1674), .IN2(\read_value_mux[7][4] ), .IN3(n1711), 
        .IN4(\read_value_mux[7][17] ), .QN(n1913) );
  OA221X1 U3082 ( .IN1(n1674), .IN2(\read_value_mux[7][4] ), .IN3(n1711), 
        .IN4(\read_value_mux[7][17] ), .IN5(n1913), .Q(n1916) );
  MUX21X1 U3083 ( .IN1(n1680), .IN2(search_data[6]), .S(\read_value_mux[7][6] ), .Q(n1915) );
  MUX21X1 U3084 ( .IN1(n1730), .IN2(search_data[27]), .S(
        \read_value_mux[7][27] ), .Q(n1914) );
  NAND4X0 U3085 ( .IN1(n1917), .IN2(n1916), .IN3(n1915), .IN4(n1914), .QN(
        n1946) );
  MUX21X1 U3086 ( .IN1(search_data[0]), .IN2(n1662), .S(\read_value_mux[7][0] ), .Q(n1924) );
  MUX21X1 U3087 ( .IN1(search_data[16]), .IN2(n1708), .S(
        \read_value_mux[7][16] ), .Q(n1923) );
  MUX21X1 U3088 ( .IN1(n1703), .IN2(search_data[14]), .S(
        \read_value_mux[7][14] ), .Q(n1921) );
  MUX21X1 U3089 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[7][24] ), .Q(n1920) );
  MUX21X1 U3090 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[7][25] ), .Q(n1919) );
  MUX21X1 U3091 ( .IN1(n1682), .IN2(search_data[7]), .S(\read_value_mux[7][7] ), .Q(n1918) );
  NAND4X0 U3092 ( .IN1(n1921), .IN2(n1920), .IN3(n1919), .IN4(n1918), .QN(
        n1922) );
  NOR4X0 U3093 ( .IN1(n1924), .IN2(n1923), .IN3(n1659), .IN4(n1922), .QN(n1944) );
  MUX21X1 U3094 ( .IN1(n1689), .IN2(search_data[9]), .S(\read_value_mux[7][9] ), .Q(n1928) );
  MUX21X1 U3095 ( .IN1(n1724), .IN2(search_data[22]), .S(
        \read_value_mux[7][22] ), .Q(n1927) );
  MUX21X1 U3096 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[7][23] ), .Q(n1926) );
  MUX21X1 U3097 ( .IN1(n1735), .IN2(search_data[29]), .S(
        \read_value_mux[7][29] ), .Q(n1925) );
  NAND4X0 U3098 ( .IN1(n1928), .IN2(n1927), .IN3(n1926), .IN4(n1925), .QN(
        n1940) );
  MUX21X1 U3099 ( .IN1(n1667), .IN2(search_data[2]), .S(\read_value_mux[7][2] ), .Q(n1932) );
  MUX21X1 U3100 ( .IN1(n1718), .IN2(search_data[20]), .S(
        \read_value_mux[7][20] ), .Q(n1931) );
  MUX21X1 U3101 ( .IN1(n1721), .IN2(search_data[21]), .S(
        \read_value_mux[7][21] ), .Q(n1930) );
  MUX21X1 U3102 ( .IN1(n1670), .IN2(search_data[3]), .S(\read_value_mux[7][3] ), .Q(n1929) );
  NAND4X0 U3103 ( .IN1(n1932), .IN2(n1931), .IN3(n1930), .IN4(n1929), .QN(
        n1939) );
  MUX21X1 U3104 ( .IN1(n1717), .IN2(search_data[19]), .S(
        \read_value_mux[7][19] ), .Q(n1936) );
  MUX21X1 U3105 ( .IN1(n1665), .IN2(search_data[1]), .S(\read_value_mux[7][1] ), .Q(n1935) );
  MUX21X1 U3106 ( .IN1(n1685), .IN2(search_data[8]), .S(\read_value_mux[7][8] ), .Q(n1934) );
  MUX21X1 U3107 ( .IN1(n1676), .IN2(search_data[5]), .S(\read_value_mux[7][5] ), .Q(n1933) );
  NAND4X0 U3108 ( .IN1(n1936), .IN2(n1935), .IN3(n1934), .IN4(n1933), .QN(
        n1937) );
  NOR4X0 U3109 ( .IN1(n1940), .IN2(n1939), .IN3(n1938), .IN4(n1937), .QN(n1943) );
  MUX21X1 U3110 ( .IN1(n1712), .IN2(search_data[18]), .S(
        \read_value_mux[7][18] ), .Q(n1941) );
  NAND4X0 U3111 ( .IN1(n1944), .IN2(n1943), .IN3(n1942), .IN4(n1941), .QN(
        n1945) );
  NOR4X0 U3112 ( .IN1(n1948), .IN2(n1947), .IN3(n1946), .IN4(n1945), .QN(n3061) );
  MUX21X1 U3113 ( .IN1(search_data[4]), .IN2(n1672), .S(\read_value_mux[6][4] ), .Q(n1957) );
  MUX21X1 U3114 ( .IN1(search_data[17]), .IN2(n1709), .S(
        \read_value_mux[6][17] ), .Q(n1956) );
  OAI22X1 U3115 ( .IN1(\read_value_mux[6][27] ), .IN2(n1732), .IN3(n1686), 
        .IN4(\read_value_mux[6][8] ), .QN(n1949) );
  AO221X1 U3116 ( .IN1(n1732), .IN2(\read_value_mux[6][27] ), .IN3(n1686), 
        .IN4(\read_value_mux[6][8] ), .IN5(n1949), .Q(n1955) );
  MUX21X1 U3117 ( .IN1(n1736), .IN2(search_data[29]), .S(
        \read_value_mux[6][29] ), .Q(n1953) );
  MUX21X1 U3118 ( .IN1(n1696), .IN2(search_data[12]), .S(
        \read_value_mux[6][12] ), .Q(n1952) );
  MUX21X1 U3119 ( .IN1(n1667), .IN2(search_data[2]), .S(\read_value_mux[6][2] ), .Q(n1951) );
  MUX21X1 U3120 ( .IN1(n1665), .IN2(search_data[1]), .S(\read_value_mux[6][1] ), .Q(n1950) );
  NAND4X0 U3121 ( .IN1(n1953), .IN2(n1952), .IN3(n1951), .IN4(n1950), .QN(
        n1954) );
  NOR4X0 U3122 ( .IN1(n1957), .IN2(n1956), .IN3(n1955), .IN4(n1954), .QN(n1989) );
  AOI22X1 U3123 ( .IN1(n1733), .IN2(\read_value_mux[6][28] ), .IN3(n1716), 
        .IN4(\read_value_mux[6][19] ), .QN(n1958) );
  OA221X1 U3124 ( .IN1(n1733), .IN2(\read_value_mux[6][28] ), .IN3(n1716), 
        .IN4(\read_value_mux[6][19] ), .IN5(n1958), .Q(n1988) );
  MUX21X1 U3125 ( .IN1(search_data[23]), .IN2(n1725), .S(
        \read_value_mux[6][23] ), .Q(n1965) );
  MUX21X1 U3126 ( .IN1(search_data[16]), .IN2(n1708), .S(
        \read_value_mux[6][16] ), .Q(n1964) );
  MUX21X1 U3127 ( .IN1(n1721), .IN2(search_data[21]), .S(
        \read_value_mux[6][21] ), .Q(n1962) );
  MUX21X1 U3128 ( .IN1(n1682), .IN2(search_data[7]), .S(\read_value_mux[6][7] ), .Q(n1961) );
  MUX21X1 U3129 ( .IN1(n1689), .IN2(search_data[9]), .S(\read_value_mux[6][9] ), .Q(n1960) );
  MUX21X1 U3130 ( .IN1(n1692), .IN2(search_data[10]), .S(
        \read_value_mux[6][10] ), .Q(n1959) );
  NAND4X0 U3131 ( .IN1(n1962), .IN2(n1961), .IN3(n1960), .IN4(n1959), .QN(
        n1963) );
  NOR4X0 U3132 ( .IN1(n1965), .IN2(n1964), .IN3(n1659), .IN4(n1963), .QN(n1987) );
  MUX21X1 U3133 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[6][24] ), .Q(n1969) );
  MUX21X1 U3134 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[6][25] ), .Q(n1968) );
  MUX21X1 U3135 ( .IN1(n1703), .IN2(search_data[14]), .S(
        \read_value_mux[6][14] ), .Q(n1967) );
  MUX21X1 U3136 ( .IN1(n1676), .IN2(search_data[5]), .S(\read_value_mux[6][5] ), .Q(n1966) );
  NAND4X0 U3137 ( .IN1(n1969), .IN2(n1968), .IN3(n1967), .IN4(n1966), .QN(
        n1985) );
  MUX21X1 U3138 ( .IN1(n1706), .IN2(n1704), .S(\read_value_mux[6][15] ), .Q(
        n1973) );
  MUX21X1 U3139 ( .IN1(n1670), .IN2(search_data[3]), .S(\read_value_mux[6][3] ), .Q(n1972) );
  MUX21X1 U3140 ( .IN1(n1739), .IN2(search_data[30]), .S(
        \read_value_mux[6][30] ), .Q(n1971) );
  MUX21X1 U3141 ( .IN1(n1712), .IN2(search_data[18]), .S(
        \read_value_mux[6][18] ), .Q(n1970) );
  NAND4X0 U3142 ( .IN1(n1973), .IN2(n1972), .IN3(n1971), .IN4(n1970), .QN(
        n1984) );
  MUX21X1 U3143 ( .IN1(n1680), .IN2(search_data[6]), .S(\read_value_mux[6][6] ), .Q(n1977) );
  MUX21X1 U3144 ( .IN1(n1724), .IN2(search_data[22]), .S(
        \read_value_mux[6][22] ), .Q(n1975) );
  MUX21X1 U3145 ( .IN1(n1695), .IN2(search_data[11]), .S(
        \read_value_mux[6][11] ), .Q(n1974) );
  NAND4X0 U3146 ( .IN1(n1977), .IN2(n1976), .IN3(n1975), .IN4(n1974), .QN(
        n1983) );
  MUX21X1 U3147 ( .IN1(n1728), .IN2(search_data[26]), .S(
        \read_value_mux[6][26] ), .Q(n1981) );
  MUX21X1 U3148 ( .IN1(n1660), .IN2(search_data[0]), .S(\read_value_mux[6][0] ), .Q(n1980) );
  MUX21X1 U3149 ( .IN1(n1718), .IN2(search_data[20]), .S(
        \read_value_mux[6][20] ), .Q(n1979) );
  MUX21X1 U3150 ( .IN1(n1741), .IN2(search_data[31]), .S(
        \read_value_mux[6][31] ), .Q(n1978) );
  NAND4X0 U3151 ( .IN1(n1981), .IN2(n1980), .IN3(n1979), .IN4(n1978), .QN(
        n1982) );
  NOR4X0 U3152 ( .IN1(n1985), .IN2(n1984), .IN3(n1983), .IN4(n1982), .QN(n1986) );
  NAND4X0 U3153 ( .IN1(n1989), .IN2(n1988), .IN3(n1987), .IN4(n1986), .QN(
        n3060) );
  MUX21X1 U3154 ( .IN1(search_data[7]), .IN2(n1681), .S(\read_value_mux[4][7] ), .Q(n1998) );
  MUX21X1 U3155 ( .IN1(search_data[11]), .IN2(n1693), .S(
        \read_value_mux[4][11] ), .Q(n1997) );
  OAI22X1 U3156 ( .IN1(n1736), .IN2(\read_value_mux[4][29] ), .IN3(n1703), 
        .IN4(\read_value_mux[4][14] ), .QN(n1990) );
  AO221X1 U3157 ( .IN1(n1736), .IN2(\read_value_mux[4][29] ), .IN3(
        \read_value_mux[4][14] ), .IN4(n1703), .IN5(n1990), .Q(n1996) );
  MUX21X1 U3158 ( .IN1(n1689), .IN2(search_data[9]), .S(\read_value_mux[4][9] ), .Q(n1994) );
  MUX21X1 U3159 ( .IN1(n1696), .IN2(search_data[12]), .S(
        \read_value_mux[4][12] ), .Q(n1993) );
  MUX21X1 U3160 ( .IN1(n1674), .IN2(search_data[4]), .S(\read_value_mux[4][4] ), .Q(n1992) );
  MUX21X1 U3161 ( .IN1(n1718), .IN2(search_data[20]), .S(
        \read_value_mux[4][20] ), .Q(n1991) );
  NAND4X0 U3162 ( .IN1(n1994), .IN2(n1993), .IN3(n1992), .IN4(n1991), .QN(
        n1995) );
  NOR4X0 U3163 ( .IN1(n1998), .IN2(n1997), .IN3(n1996), .IN4(n1995), .QN(n2030) );
  AOI22X1 U3164 ( .IN1(n1668), .IN2(\read_value_mux[4][2] ), .IN3(n1724), 
        .IN4(\read_value_mux[4][22] ), .QN(n1999) );
  OA221X1 U3165 ( .IN1(n1668), .IN2(\read_value_mux[4][2] ), .IN3(n1724), 
        .IN4(\read_value_mux[4][22] ), .IN5(n1999), .Q(n2029) );
  MUX21X1 U3166 ( .IN1(search_data[23]), .IN2(n1725), .S(
        \read_value_mux[4][23] ), .Q(n2006) );
  MUX21X1 U3167 ( .IN1(search_data[31]), .IN2(n1740), .S(
        \read_value_mux[4][31] ), .Q(n2005) );
  MUX21X1 U3168 ( .IN1(n1716), .IN2(search_data[19]), .S(
        \read_value_mux[4][19] ), .Q(n2003) );
  MUX21X1 U3169 ( .IN1(n1670), .IN2(search_data[3]), .S(\read_value_mux[4][3] ), .Q(n2002) );
  MUX21X1 U3170 ( .IN1(n1676), .IN2(search_data[5]), .S(\read_value_mux[4][5] ), .Q(n2001) );
  NAND4X0 U3171 ( .IN1(n2003), .IN2(n2002), .IN3(n2001), .IN4(n2000), .QN(
        n2004) );
  NOR4X0 U3172 ( .IN1(n2006), .IN2(n2005), .IN3(n1659), .IN4(n2004), .QN(n2028) );
  MUX21X1 U3173 ( .IN1(n1711), .IN2(search_data[17]), .S(
        \read_value_mux[4][17] ), .Q(n2010) );
  MUX21X1 U3174 ( .IN1(n1738), .IN2(search_data[30]), .S(
        \read_value_mux[4][30] ), .Q(n2009) );
  MUX21X1 U3175 ( .IN1(n1660), .IN2(search_data[0]), .S(\read_value_mux[4][0] ), .Q(n2008) );
  NAND4X0 U3176 ( .IN1(n2010), .IN2(n2009), .IN3(n2008), .IN4(n2007), .QN(
        n2026) );
  MUX21X1 U3177 ( .IN1(n1714), .IN2(search_data[18]), .S(
        \read_value_mux[4][18] ), .Q(n2014) );
  MUX21X1 U3178 ( .IN1(n1708), .IN2(search_data[16]), .S(
        \read_value_mux[4][16] ), .Q(n2013) );
  MUX21X1 U3179 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[4][25] ), .Q(n2012) );
  MUX21X1 U3180 ( .IN1(n1705), .IN2(n1704), .S(\read_value_mux[4][15] ), .Q(
        n2011) );
  NAND4X0 U3181 ( .IN1(n2014), .IN2(n2013), .IN3(n2012), .IN4(n2011), .QN(
        n2025) );
  MUX21X1 U3182 ( .IN1(n1685), .IN2(search_data[8]), .S(\read_value_mux[4][8] ), .Q(n2018) );
  MUX21X1 U3183 ( .IN1(n1720), .IN2(search_data[21]), .S(
        \read_value_mux[4][21] ), .Q(n2017) );
  MUX21X1 U3184 ( .IN1(n1665), .IN2(search_data[1]), .S(\read_value_mux[4][1] ), .Q(n2016) );
  MUX21X1 U3185 ( .IN1(n1680), .IN2(search_data[6]), .S(\read_value_mux[4][6] ), .Q(n2015) );
  NAND4X0 U3186 ( .IN1(n2018), .IN2(n2017), .IN3(n2016), .IN4(n2015), .QN(
        n2024) );
  MUX21X1 U3187 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[4][24] ), .Q(n2022) );
  MUX21X1 U3188 ( .IN1(n1691), .IN2(n1690), .S(\read_value_mux[4][10] ), .Q(
        n2021) );
  MUX21X1 U3189 ( .IN1(n1730), .IN2(search_data[27]), .S(
        \read_value_mux[4][27] ), .Q(n2020) );
  MUX21X1 U3190 ( .IN1(n1728), .IN2(search_data[26]), .S(
        \read_value_mux[4][26] ), .Q(n2019) );
  NAND4X0 U3191 ( .IN1(n2022), .IN2(n2021), .IN3(n2020), .IN4(n2019), .QN(
        n2023) );
  NOR4X0 U3192 ( .IN1(n2026), .IN2(n2025), .IN3(n2024), .IN4(n2023), .QN(n2027) );
  NAND4X0 U3193 ( .IN1(n2030), .IN2(n2029), .IN3(n2028), .IN4(n2027), .QN(
        n3057) );
  MUX21X1 U3194 ( .IN1(search_data[29]), .IN2(n1734), .S(
        \read_value_mux[1][29] ), .Q(n2071) );
  MUX21X1 U3195 ( .IN1(n1690), .IN2(n1691), .S(\read_value_mux[1][10] ), .Q(
        n2070) );
  AOI22X1 U3196 ( .IN1(n1727), .IN2(\read_value_mux[1][25] ), .IN3(n1716), 
        .IN4(\read_value_mux[1][19] ), .QN(n2031) );
  OA221X1 U3197 ( .IN1(n1727), .IN2(\read_value_mux[1][25] ), .IN3(n1717), 
        .IN4(\read_value_mux[1][19] ), .IN5(n2031), .Q(n2036) );
  AOI22X1 U3198 ( .IN1(n1677), .IN2(\read_value_mux[1][5] ), .IN3(n1671), 
        .IN4(\read_value_mux[1][3] ), .QN(n2032) );
  OA221X1 U3199 ( .IN1(n1677), .IN2(\read_value_mux[1][5] ), .IN3(n1671), 
        .IN4(\read_value_mux[1][3] ), .IN5(n2032), .Q(n2035) );
  MUX21X1 U3200 ( .IN1(n1728), .IN2(search_data[26]), .S(
        \read_value_mux[1][26] ), .Q(n2034) );
  MUX21X1 U3201 ( .IN1(n1705), .IN2(n1704), .S(\read_value_mux[1][15] ), .Q(
        n2033) );
  NAND4X0 U3202 ( .IN1(n2036), .IN2(n2035), .IN3(n2034), .IN4(n2033), .QN(
        n2069) );
  MUX21X1 U3203 ( .IN1(search_data[20]), .IN2(n1718), .S(
        \read_value_mux[1][20] ), .Q(n2043) );
  MUX21X1 U3204 ( .IN1(search_data[7]), .IN2(n1681), .S(\read_value_mux[1][7] ), .Q(n2042) );
  MUX21X1 U3205 ( .IN1(n1720), .IN2(search_data[21]), .S(
        \read_value_mux[1][21] ), .Q(n2040) );
  MUX21X1 U3206 ( .IN1(n1702), .IN2(search_data[14]), .S(
        \read_value_mux[1][14] ), .Q(n2039) );
  MUX21X1 U3207 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[1][24] ), .Q(n2038) );
  MUX21X1 U3208 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[1][28] ), .Q(n2037) );
  NAND4X0 U3209 ( .IN1(n2040), .IN2(n2039), .IN3(n2038), .IN4(n2037), .QN(
        n2041) );
  NOR4X0 U3210 ( .IN1(n2043), .IN2(n2042), .IN3(n1659), .IN4(n2041), .QN(n2067) );
  MUX21X1 U3211 ( .IN1(n1699), .IN2(search_data[13]), .S(
        \read_value_mux[1][13] ), .Q(n2047) );
  MUX21X1 U3212 ( .IN1(n1667), .IN2(search_data[2]), .S(\read_value_mux[1][2] ), .Q(n2046) );
  MUX21X1 U3213 ( .IN1(n1661), .IN2(search_data[0]), .S(\read_value_mux[1][0] ), .Q(n2045) );
  MUX21X1 U3214 ( .IN1(n1723), .IN2(search_data[22]), .S(
        \read_value_mux[1][22] ), .Q(n2044) );
  NAND4X0 U3215 ( .IN1(n2047), .IN2(n2046), .IN3(n2045), .IN4(n2044), .QN(
        n2063) );
  MUX21X1 U3216 ( .IN1(n1679), .IN2(search_data[6]), .S(\read_value_mux[1][6] ), .Q(n2051) );
  MUX21X1 U3217 ( .IN1(n1707), .IN2(search_data[16]), .S(
        \read_value_mux[1][16] ), .Q(n2050) );
  MUX21X1 U3218 ( .IN1(n1695), .IN2(search_data[11]), .S(
        \read_value_mux[1][11] ), .Q(n2049) );
  MUX21X1 U3219 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[1][23] ), .Q(n2048) );
  NAND4X0 U3220 ( .IN1(n2051), .IN2(n2050), .IN3(n2049), .IN4(n2048), .QN(
        n2062) );
  MUX21X1 U3221 ( .IN1(n1710), .IN2(search_data[17]), .S(
        \read_value_mux[1][17] ), .Q(n2055) );
  MUX21X1 U3222 ( .IN1(n1738), .IN2(search_data[30]), .S(
        \read_value_mux[1][30] ), .Q(n2054) );
  MUX21X1 U3223 ( .IN1(n1730), .IN2(search_data[27]), .S(
        \read_value_mux[1][27] ), .Q(n2053) );
  MUX21X1 U3224 ( .IN1(n1664), .IN2(search_data[1]), .S(\read_value_mux[1][1] ), .Q(n2052) );
  NAND4X0 U3225 ( .IN1(n2055), .IN2(n2054), .IN3(n2053), .IN4(n2052), .QN(
        n2061) );
  MUX21X1 U3226 ( .IN1(n1696), .IN2(search_data[12]), .S(
        \read_value_mux[1][12] ), .Q(n2059) );
  MUX21X1 U3227 ( .IN1(n1685), .IN2(search_data[8]), .S(\read_value_mux[1][8] ), .Q(n2058) );
  MUX21X1 U3228 ( .IN1(n1713), .IN2(search_data[18]), .S(
        \read_value_mux[1][18] ), .Q(n2057) );
  MUX21X1 U3229 ( .IN1(n1741), .IN2(search_data[31]), .S(
        \read_value_mux[1][31] ), .Q(n2056) );
  NAND4X0 U3230 ( .IN1(n2059), .IN2(n2058), .IN3(n2057), .IN4(n2056), .QN(
        n2060) );
  NOR4X0 U3231 ( .IN1(n2063), .IN2(n2062), .IN3(n2061), .IN4(n2060), .QN(n2066) );
  MUX21X1 U3232 ( .IN1(n1673), .IN2(search_data[4]), .S(\read_value_mux[1][4] ), .Q(n2065) );
  MUX21X1 U3233 ( .IN1(n1688), .IN2(search_data[9]), .S(\read_value_mux[1][9] ), .Q(n2064) );
  NAND4X0 U3234 ( .IN1(n2067), .IN2(n2066), .IN3(n2065), .IN4(n2064), .QN(
        n2068) );
  NOR4X0 U3235 ( .IN1(n2071), .IN2(n2070), .IN3(n2069), .IN4(n2068), .QN(n3118) );
  MUX21X1 U3236 ( .IN1(search_data[19]), .IN2(n1715), .S(
        \read_value_mux[9][19] ), .Q(n2080) );
  MUX21X1 U3237 ( .IN1(search_data[18]), .IN2(n1714), .S(
        \read_value_mux[9][18] ), .Q(n2079) );
  OAI22X1 U3238 ( .IN1(n1718), .IN2(\read_value_mux[9][20] ), .IN3(n1711), 
        .IN4(\read_value_mux[9][17] ), .QN(n2072) );
  AO221X1 U3239 ( .IN1(n1718), .IN2(\read_value_mux[9][20] ), .IN3(
        \read_value_mux[9][17] ), .IN4(n1711), .IN5(n2072), .Q(n2078) );
  MUX21X1 U3240 ( .IN1(n1699), .IN2(search_data[13]), .S(
        \read_value_mux[9][13] ), .Q(n2076) );
  MUX21X1 U3241 ( .IN1(n1705), .IN2(n1704), .S(\read_value_mux[9][15] ), .Q(
        n2075) );
  MUX21X1 U3242 ( .IN1(n1730), .IN2(search_data[27]), .S(
        \read_value_mux[9][27] ), .Q(n2074) );
  MUX21X1 U3243 ( .IN1(n1679), .IN2(search_data[6]), .S(\read_value_mux[9][6] ), .Q(n2073) );
  NAND4X0 U3244 ( .IN1(n2076), .IN2(n2075), .IN3(n2074), .IN4(n2073), .QN(
        n2077) );
  NOR4X0 U3245 ( .IN1(n2080), .IN2(n2079), .IN3(n2078), .IN4(n2077), .QN(n2112) );
  AOI22X1 U3246 ( .IN1(n1683), .IN2(\read_value_mux[9][7] ), .IN3(n1697), 
        .IN4(\read_value_mux[9][12] ), .QN(n2081) );
  OA221X1 U3247 ( .IN1(n1683), .IN2(\read_value_mux[9][7] ), .IN3(n1697), 
        .IN4(\read_value_mux[9][12] ), .IN5(n2081), .Q(n2111) );
  MUX21X1 U3248 ( .IN1(search_data[4]), .IN2(n1672), .S(\read_value_mux[9][4] ), .Q(n2088) );
  MUX21X1 U3249 ( .IN1(search_data[29]), .IN2(n1734), .S(
        \read_value_mux[9][29] ), .Q(n2087) );
  MUX21X1 U3250 ( .IN1(n1662), .IN2(search_data[0]), .S(\read_value_mux[9][0] ), .Q(n2085) );
  MUX21X1 U3251 ( .IN1(n1689), .IN2(search_data[9]), .S(\read_value_mux[9][9] ), .Q(n2084) );
  MUX21X1 U3252 ( .IN1(n1723), .IN2(search_data[22]), .S(
        \read_value_mux[9][22] ), .Q(n2083) );
  MUX21X1 U3253 ( .IN1(n1667), .IN2(search_data[2]), .S(\read_value_mux[9][2] ), .Q(n2082) );
  NAND4X0 U3254 ( .IN1(n2085), .IN2(n2084), .IN3(n2083), .IN4(n2082), .QN(
        n2086) );
  NOR4X0 U3255 ( .IN1(n2088), .IN2(n2087), .IN3(n1659), .IN4(n2086), .QN(n2110) );
  MUX21X1 U3256 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[9][24] ), .Q(n2092) );
  MUX21X1 U3257 ( .IN1(n1670), .IN2(search_data[3]), .S(\read_value_mux[9][3] ), .Q(n2091) );
  MUX21X1 U3258 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[9][25] ), .Q(n2090) );
  MUX21X1 U3259 ( .IN1(n1741), .IN2(search_data[31]), .S(
        \read_value_mux[9][31] ), .Q(n2089) );
  NAND4X0 U3260 ( .IN1(n2092), .IN2(n2091), .IN3(n2090), .IN4(n2089), .QN(
        n2108) );
  MUX21X1 U3261 ( .IN1(n1729), .IN2(search_data[26]), .S(
        \read_value_mux[9][26] ), .Q(n2096) );
  MUX21X1 U3262 ( .IN1(n1694), .IN2(search_data[11]), .S(
        \read_value_mux[9][11] ), .Q(n2095) );
  MUX21X1 U3263 ( .IN1(n1685), .IN2(search_data[8]), .S(\read_value_mux[9][8] ), .Q(n2094) );
  MUX21X1 U3264 ( .IN1(n1707), .IN2(search_data[16]), .S(
        \read_value_mux[9][16] ), .Q(n2093) );
  NAND4X0 U3265 ( .IN1(n2096), .IN2(n2095), .IN3(n2094), .IN4(n2093), .QN(
        n2107) );
  MUX21X1 U3266 ( .IN1(n1702), .IN2(search_data[14]), .S(
        \read_value_mux[9][14] ), .Q(n2100) );
  MUX21X1 U3267 ( .IN1(n1676), .IN2(search_data[5]), .S(\read_value_mux[9][5] ), .Q(n2099) );
  MUX21X1 U3268 ( .IN1(n1691), .IN2(n1690), .S(\read_value_mux[9][10] ), .Q(
        n2098) );
  NAND4X0 U3269 ( .IN1(n2100), .IN2(n2099), .IN3(n2098), .IN4(n2097), .QN(
        n2106) );
  MUX21X1 U3270 ( .IN1(n1664), .IN2(search_data[1]), .S(\read_value_mux[9][1] ), .Q(n2104) );
  MUX21X1 U3271 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[9][23] ), .Q(n2103) );
  MUX21X1 U3272 ( .IN1(n1738), .IN2(search_data[30]), .S(
        \read_value_mux[9][30] ), .Q(n2102) );
  MUX21X1 U3273 ( .IN1(n1720), .IN2(search_data[21]), .S(
        \read_value_mux[9][21] ), .Q(n2101) );
  NAND4X0 U3274 ( .IN1(n2104), .IN2(n2103), .IN3(n2102), .IN4(n2101), .QN(
        n2105) );
  NOR4X0 U3275 ( .IN1(n2108), .IN2(n2107), .IN3(n2106), .IN4(n2105), .QN(n2109) );
  NAND4X0 U3276 ( .IN1(n2112), .IN2(n2111), .IN3(n2110), .IN4(n2109), .QN(
        n3094) );
  MUX21X1 U3277 ( .IN1(search_data[28]), .IN2(n1733), .S(
        \read_value_mux[10][28] ), .Q(n2153) );
  MUX21X1 U3278 ( .IN1(n1704), .IN2(n1705), .S(\read_value_mux[10][15] ), .Q(
        n2152) );
  AOI22X1 U3279 ( .IN1(n1661), .IN2(\read_value_mux[10][0] ), .IN3(n1736), 
        .IN4(\read_value_mux[10][29] ), .QN(n2113) );
  OA221X1 U3280 ( .IN1(n1661), .IN2(\read_value_mux[10][0] ), .IN3(n1736), 
        .IN4(\read_value_mux[10][29] ), .IN5(n2113), .Q(n2118) );
  AOI22X1 U3281 ( .IN1(n1691), .IN2(\read_value_mux[10][10] ), .IN3(n1671), 
        .IN4(\read_value_mux[10][3] ), .QN(n2114) );
  OA221X1 U3282 ( .IN1(n1691), .IN2(\read_value_mux[10][10] ), .IN3(n1671), 
        .IN4(\read_value_mux[10][3] ), .IN5(n2114), .Q(n2117) );
  MUX21X1 U3283 ( .IN1(n1694), .IN2(search_data[11]), .S(
        \read_value_mux[10][11] ), .Q(n2116) );
  MUX21X1 U3284 ( .IN1(n1738), .IN2(search_data[30]), .S(
        \read_value_mux[10][30] ), .Q(n2115) );
  NAND4X0 U3285 ( .IN1(n2118), .IN2(n2117), .IN3(n2116), .IN4(n2115), .QN(
        n2151) );
  MUX21X1 U3286 ( .IN1(search_data[14]), .IN2(n1701), .S(
        \read_value_mux[10][14] ), .Q(n2125) );
  MUX21X1 U3287 ( .IN1(search_data[26]), .IN2(n1728), .S(
        \read_value_mux[10][26] ), .Q(n2124) );
  MUX21X1 U3288 ( .IN1(n1685), .IN2(search_data[8]), .S(
        \read_value_mux[10][8] ), .Q(n2122) );
  MUX21X1 U3289 ( .IN1(n1723), .IN2(search_data[22]), .S(
        \read_value_mux[10][22] ), .Q(n2121) );
  MUX21X1 U3290 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[10][25] ), .Q(n2120) );
  MUX21X1 U3291 ( .IN1(n1696), .IN2(search_data[12]), .S(
        \read_value_mux[10][12] ), .Q(n2119) );
  NAND4X0 U3292 ( .IN1(n2122), .IN2(n2121), .IN3(n2120), .IN4(n2119), .QN(
        n2123) );
  NOR4X0 U3293 ( .IN1(n2125), .IN2(n2124), .IN3(n1659), .IN4(n2123), .QN(n2149) );
  MUX21X1 U3294 ( .IN1(n1673), .IN2(search_data[4]), .S(
        \read_value_mux[10][4] ), .Q(n2129) );
  MUX21X1 U3295 ( .IN1(n1688), .IN2(search_data[9]), .S(
        \read_value_mux[10][9] ), .Q(n2128) );
  MUX21X1 U3296 ( .IN1(n1679), .IN2(search_data[6]), .S(
        \read_value_mux[10][6] ), .Q(n2127) );
  MUX21X1 U3297 ( .IN1(n1710), .IN2(search_data[17]), .S(
        \read_value_mux[10][17] ), .Q(n2126) );
  NAND4X0 U3298 ( .IN1(n2129), .IN2(n2128), .IN3(n2127), .IN4(n2126), .QN(
        n2145) );
  MUX21X1 U3299 ( .IN1(n1713), .IN2(search_data[18]), .S(
        \read_value_mux[10][18] ), .Q(n2133) );
  MUX21X1 U3300 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[10][24] ), .Q(n2132) );
  MUX21X1 U3301 ( .IN1(n1740), .IN2(search_data[31]), .S(
        \read_value_mux[10][31] ), .Q(n2131) );
  MUX21X1 U3302 ( .IN1(n1664), .IN2(search_data[1]), .S(
        \read_value_mux[10][1] ), .Q(n2130) );
  NAND4X0 U3303 ( .IN1(n2133), .IN2(n2132), .IN3(n2131), .IN4(n2130), .QN(
        n2144) );
  MUX21X1 U3304 ( .IN1(n1718), .IN2(search_data[20]), .S(
        \read_value_mux[10][20] ), .Q(n2137) );
  MUX21X1 U3305 ( .IN1(n1682), .IN2(search_data[7]), .S(
        \read_value_mux[10][7] ), .Q(n2136) );
  MUX21X1 U3306 ( .IN1(n1667), .IN2(search_data[2]), .S(
        \read_value_mux[10][2] ), .Q(n2135) );
  MUX21X1 U3307 ( .IN1(n1720), .IN2(search_data[21]), .S(
        \read_value_mux[10][21] ), .Q(n2134) );
  NAND4X0 U3308 ( .IN1(n2137), .IN2(n2136), .IN3(n2135), .IN4(n2134), .QN(
        n2143) );
  MUX21X1 U3309 ( .IN1(n1676), .IN2(search_data[5]), .S(
        \read_value_mux[10][5] ), .Q(n2141) );
  MUX21X1 U3310 ( .IN1(n1731), .IN2(search_data[27]), .S(
        \read_value_mux[10][27] ), .Q(n2140) );
  MUX21X1 U3311 ( .IN1(n1699), .IN2(search_data[13]), .S(
        \read_value_mux[10][13] ), .Q(n2139) );
  MUX21X1 U3312 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[10][23] ), .Q(n2138) );
  NAND4X0 U3313 ( .IN1(n2141), .IN2(n2140), .IN3(n2139), .IN4(n2138), .QN(
        n2142) );
  NOR4X0 U3314 ( .IN1(n2145), .IN2(n2144), .IN3(n2143), .IN4(n2142), .QN(n2148) );
  MUX21X1 U3315 ( .IN1(n1715), .IN2(search_data[19]), .S(
        \read_value_mux[10][19] ), .Q(n2147) );
  MUX21X1 U3316 ( .IN1(n1707), .IN2(search_data[16]), .S(
        \read_value_mux[10][16] ), .Q(n2146) );
  NAND4X0 U3317 ( .IN1(n2149), .IN2(n2148), .IN3(n2147), .IN4(n2146), .QN(
        n2150) );
  NOR4X0 U3318 ( .IN1(n2153), .IN2(n2152), .IN3(n2151), .IN4(n2150), .QN(n3064) );
  OAI22X1 U3319 ( .IN1(\read_value_mux[16][5] ), .IN2(n1677), .IN3(n1683), 
        .IN4(\read_value_mux[16][7] ), .QN(n2154) );
  AO221X1 U3320 ( .IN1(n1676), .IN2(\read_value_mux[16][5] ), .IN3(n1683), 
        .IN4(\read_value_mux[16][7] ), .IN5(n2154), .Q(n2194) );
  OAI22X1 U3321 ( .IN1(\read_value_mux[16][29] ), .IN2(n1736), .IN3(n1668), 
        .IN4(\read_value_mux[16][2] ), .QN(n2155) );
  AO221X1 U3322 ( .IN1(n1736), .IN2(\read_value_mux[16][29] ), .IN3(n1668), 
        .IN4(\read_value_mux[16][2] ), .IN5(n2155), .Q(n2193) );
  MUX21X1 U3323 ( .IN1(n1660), .IN2(search_data[0]), .S(
        \read_value_mux[16][0] ), .Q(n2159) );
  MUX21X1 U3324 ( .IN1(n1723), .IN2(search_data[22]), .S(
        \read_value_mux[16][22] ), .Q(n2158) );
  MUX21X1 U3325 ( .IN1(n1688), .IN2(search_data[9]), .S(
        \read_value_mux[16][9] ), .Q(n2157) );
  MUX21X1 U3326 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[16][25] ), .Q(n2156) );
  NAND4X0 U3327 ( .IN1(n2159), .IN2(n2158), .IN3(n2157), .IN4(n2156), .QN(
        n2192) );
  MUX21X1 U3328 ( .IN1(search_data[16]), .IN2(n1708), .S(
        \read_value_mux[16][16] ), .Q(n2166) );
  MUX21X1 U3329 ( .IN1(search_data[28]), .IN2(n1733), .S(
        \read_value_mux[16][28] ), .Q(n2165) );
  MUX21X1 U3330 ( .IN1(n1679), .IN2(search_data[6]), .S(
        \read_value_mux[16][6] ), .Q(n2163) );
  MUX21X1 U3331 ( .IN1(n1738), .IN2(search_data[30]), .S(
        \read_value_mux[16][30] ), .Q(n2162) );
  MUX21X1 U3332 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[16][24] ), .Q(n2161) );
  MUX21X1 U3333 ( .IN1(n1673), .IN2(search_data[4]), .S(
        \read_value_mux[16][4] ), .Q(n2160) );
  NAND4X0 U3334 ( .IN1(n2163), .IN2(n2162), .IN3(n2161), .IN4(n2160), .QN(
        n2164) );
  NOR4X0 U3335 ( .IN1(n2166), .IN2(n2165), .IN3(n1659), .IN4(n2164), .QN(n2190) );
  MUX21X1 U3336 ( .IN1(n1705), .IN2(n1704), .S(\read_value_mux[16][15] ), .Q(
        n2170) );
  MUX21X1 U3337 ( .IN1(n1741), .IN2(search_data[31]), .S(
        \read_value_mux[16][31] ), .Q(n2169) );
  MUX21X1 U3338 ( .IN1(n1718), .IN2(search_data[20]), .S(
        \read_value_mux[16][20] ), .Q(n2168) );
  MUX21X1 U3339 ( .IN1(n1710), .IN2(search_data[17]), .S(
        \read_value_mux[16][17] ), .Q(n2167) );
  NAND4X0 U3340 ( .IN1(n2170), .IN2(n2169), .IN3(n2168), .IN4(n2167), .QN(
        n2186) );
  MUX21X1 U3341 ( .IN1(n1692), .IN2(n1690), .S(\read_value_mux[16][10] ), .Q(
        n2174) );
  MUX21X1 U3342 ( .IN1(n1716), .IN2(search_data[19]), .S(
        \read_value_mux[16][19] ), .Q(n2173) );
  MUX21X1 U3343 ( .IN1(n1664), .IN2(search_data[1]), .S(
        \read_value_mux[16][1] ), .Q(n2172) );
  MUX21X1 U3344 ( .IN1(n1685), .IN2(search_data[8]), .S(
        \read_value_mux[16][8] ), .Q(n2171) );
  NAND4X0 U3345 ( .IN1(n2174), .IN2(n2173), .IN3(n2172), .IN4(n2171), .QN(
        n2185) );
  MUX21X1 U3346 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[16][23] ), .Q(n2178) );
  MUX21X1 U3347 ( .IN1(n1713), .IN2(search_data[18]), .S(
        \read_value_mux[16][18] ), .Q(n2177) );
  MUX21X1 U3348 ( .IN1(n1696), .IN2(search_data[12]), .S(
        \read_value_mux[16][12] ), .Q(n2176) );
  MUX21X1 U3349 ( .IN1(n1702), .IN2(search_data[14]), .S(
        \read_value_mux[16][14] ), .Q(n2175) );
  NAND4X0 U3350 ( .IN1(n2178), .IN2(n2177), .IN3(n2176), .IN4(n2175), .QN(
        n2184) );
  MUX21X1 U3351 ( .IN1(n1720), .IN2(search_data[21]), .S(
        \read_value_mux[16][21] ), .Q(n2182) );
  MUX21X1 U3352 ( .IN1(n1731), .IN2(search_data[27]), .S(
        \read_value_mux[16][27] ), .Q(n2181) );
  MUX21X1 U3353 ( .IN1(n1670), .IN2(search_data[3]), .S(
        \read_value_mux[16][3] ), .Q(n2180) );
  MUX21X1 U3354 ( .IN1(n1694), .IN2(search_data[11]), .S(
        \read_value_mux[16][11] ), .Q(n2179) );
  NAND4X0 U3355 ( .IN1(n2182), .IN2(n2181), .IN3(n2180), .IN4(n2179), .QN(
        n2183) );
  NOR4X0 U3356 ( .IN1(n2186), .IN2(n2185), .IN3(n2184), .IN4(n2183), .QN(n2189) );
  MUX21X1 U3357 ( .IN1(n1729), .IN2(search_data[26]), .S(
        \read_value_mux[16][26] ), .Q(n2188) );
  MUX21X1 U3358 ( .IN1(n1699), .IN2(search_data[13]), .S(
        \read_value_mux[16][13] ), .Q(n2187) );
  NAND4X0 U3359 ( .IN1(n2190), .IN2(n2189), .IN3(n2188), .IN4(n2187), .QN(
        n2191) );
  NOR4X0 U3360 ( .IN1(n2194), .IN2(n2193), .IN3(n2192), .IN4(n2191), .QN(n3087) );
  MUX21X1 U3361 ( .IN1(search_data[14]), .IN2(n1701), .S(
        \read_value_mux[14][14] ), .Q(n2203) );
  MUX21X1 U3362 ( .IN1(search_data[28]), .IN2(n1733), .S(
        \read_value_mux[14][28] ), .Q(n2202) );
  OAI22X1 U3363 ( .IN1(n1708), .IN2(\read_value_mux[14][16] ), .IN3(n1668), 
        .IN4(\read_value_mux[14][2] ), .QN(n2195) );
  AO221X1 U3364 ( .IN1(n1708), .IN2(\read_value_mux[14][16] ), .IN3(
        \read_value_mux[14][2] ), .IN4(n1668), .IN5(n2195), .Q(n2201) );
  MUX21X1 U3365 ( .IN1(n1741), .IN2(search_data[31]), .S(
        \read_value_mux[14][31] ), .Q(n2199) );
  MUX21X1 U3366 ( .IN1(n1661), .IN2(search_data[0]), .S(
        \read_value_mux[14][0] ), .Q(n2198) );
  MUX21X1 U3367 ( .IN1(n1699), .IN2(search_data[13]), .S(
        \read_value_mux[14][13] ), .Q(n2197) );
  MUX21X1 U3368 ( .IN1(n1676), .IN2(search_data[5]), .S(
        \read_value_mux[14][5] ), .Q(n2196) );
  NAND4X0 U3369 ( .IN1(n2199), .IN2(n2198), .IN3(n2197), .IN4(n2196), .QN(
        n2200) );
  NOR4X0 U3370 ( .IN1(n2203), .IN2(n2202), .IN3(n2201), .IN4(n2200), .QN(n2235) );
  AOI22X1 U3371 ( .IN1(n1725), .IN2(\read_value_mux[14][23] ), .IN3(n1706), 
        .IN4(\read_value_mux[14][15] ), .QN(n2204) );
  OA221X1 U3372 ( .IN1(n1725), .IN2(\read_value_mux[14][23] ), .IN3(n1706), 
        .IN4(\read_value_mux[14][15] ), .IN5(n2204), .Q(n2234) );
  MUX21X1 U3373 ( .IN1(search_data[11]), .IN2(n1693), .S(
        \read_value_mux[14][11] ), .Q(n2211) );
  MUX21X1 U3374 ( .IN1(search_data[21]), .IN2(n1719), .S(
        \read_value_mux[14][21] ), .Q(n2210) );
  MUX21X1 U3375 ( .IN1(n1670), .IN2(search_data[3]), .S(
        \read_value_mux[14][3] ), .Q(n2208) );
  MUX21X1 U3376 ( .IN1(n1685), .IN2(search_data[8]), .S(
        \read_value_mux[14][8] ), .Q(n2207) );
  MUX21X1 U3377 ( .IN1(n1664), .IN2(search_data[1]), .S(
        \read_value_mux[14][1] ), .Q(n2206) );
  MUX21X1 U3378 ( .IN1(n1738), .IN2(search_data[30]), .S(
        \read_value_mux[14][30] ), .Q(n2205) );
  NAND4X0 U3379 ( .IN1(n2208), .IN2(n2207), .IN3(n2206), .IN4(n2205), .QN(
        n2209) );
  NOR4X0 U3380 ( .IN1(n2211), .IN2(n2210), .IN3(n1659), .IN4(n2209), .QN(n2233) );
  MUX21X1 U3381 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[14][25] ), .Q(n2215) );
  MUX21X1 U3382 ( .IN1(n1696), .IN2(search_data[12]), .S(
        \read_value_mux[14][12] ), .Q(n2214) );
  MUX21X1 U3383 ( .IN1(n1713), .IN2(search_data[18]), .S(
        \read_value_mux[14][18] ), .Q(n2213) );
  MUX21X1 U3384 ( .IN1(n1729), .IN2(search_data[26]), .S(
        \read_value_mux[14][26] ), .Q(n2212) );
  NAND4X0 U3385 ( .IN1(n2215), .IN2(n2214), .IN3(n2213), .IN4(n2212), .QN(
        n2231) );
  MUX21X1 U3386 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[14][24] ), .Q(n2219) );
  MUX21X1 U3387 ( .IN1(n1679), .IN2(search_data[6]), .S(
        \read_value_mux[14][6] ), .Q(n2218) );
  MUX21X1 U3388 ( .IN1(n1710), .IN2(search_data[17]), .S(
        \read_value_mux[14][17] ), .Q(n2217) );
  MUX21X1 U3389 ( .IN1(n1716), .IN2(search_data[19]), .S(
        \read_value_mux[14][19] ), .Q(n2216) );
  NAND4X0 U3390 ( .IN1(n2219), .IN2(n2218), .IN3(n2217), .IN4(n2216), .QN(
        n2230) );
  MUX21X1 U3391 ( .IN1(n1682), .IN2(search_data[7]), .S(
        \read_value_mux[14][7] ), .Q(n2223) );
  MUX21X1 U3392 ( .IN1(n1730), .IN2(search_data[27]), .S(
        \read_value_mux[14][27] ), .Q(n2222) );
  MUX21X1 U3393 ( .IN1(n1692), .IN2(n1690), .S(\read_value_mux[14][10] ), .Q(
        n2221) );
  MUX21X1 U3394 ( .IN1(n1718), .IN2(search_data[20]), .S(
        \read_value_mux[14][20] ), .Q(n2220) );
  NAND4X0 U3395 ( .IN1(n2223), .IN2(n2222), .IN3(n2221), .IN4(n2220), .QN(
        n2229) );
  MUX21X1 U3396 ( .IN1(n1688), .IN2(search_data[9]), .S(
        \read_value_mux[14][9] ), .Q(n2227) );
  MUX21X1 U3397 ( .IN1(n1723), .IN2(search_data[22]), .S(
        \read_value_mux[14][22] ), .Q(n2226) );
  MUX21X1 U3398 ( .IN1(n1673), .IN2(search_data[4]), .S(
        \read_value_mux[14][4] ), .Q(n2225) );
  MUX21X1 U3399 ( .IN1(n1735), .IN2(search_data[29]), .S(
        \read_value_mux[14][29] ), .Q(n2224) );
  NAND4X0 U3400 ( .IN1(n2227), .IN2(n2226), .IN3(n2225), .IN4(n2224), .QN(
        n2228) );
  NOR4X0 U3401 ( .IN1(n2231), .IN2(n2230), .IN3(n2229), .IN4(n2228), .QN(n2232) );
  NAND4X0 U3402 ( .IN1(n2235), .IN2(n2234), .IN3(n2233), .IN4(n2232), .QN(
        n3088) );
  MUX21X1 U3403 ( .IN1(search_data[11]), .IN2(n1693), .S(
        \read_value_mux[12][11] ), .Q(n2240) );
  MUX21X1 U3404 ( .IN1(search_data[2]), .IN2(n1666), .S(
        \read_value_mux[12][2] ), .Q(n2239) );
  OAI22X1 U3405 ( .IN1(\read_value_mux[12][30] ), .IN2(n1739), .IN3(n1708), 
        .IN4(\read_value_mux[12][16] ), .QN(n2236) );
  AO221X1 U3406 ( .IN1(n1739), .IN2(\read_value_mux[12][30] ), .IN3(n1708), 
        .IN4(\read_value_mux[12][16] ), .IN5(n2236), .Q(n2238) );
  NOR4X0 U3407 ( .IN1(n2240), .IN2(n2239), .IN3(n2238), .IN4(n2237), .QN(n2272) );
  AOI22X1 U3408 ( .IN1(n1683), .IN2(\read_value_mux[12][7] ), .IN3(n1728), 
        .IN4(\read_value_mux[12][26] ), .QN(n2241) );
  OA221X1 U3409 ( .IN1(n1683), .IN2(\read_value_mux[12][7] ), .IN3(n1728), 
        .IN4(\read_value_mux[12][26] ), .IN5(n2241), .Q(n2271) );
  MUX21X1 U3410 ( .IN1(search_data[10]), .IN2(n1691), .S(
        \read_value_mux[12][10] ), .Q(n2248) );
  MUX21X1 U3411 ( .IN1(search_data[6]), .IN2(n1678), .S(
        \read_value_mux[12][6] ), .Q(n2247) );
  MUX21X1 U3412 ( .IN1(n1720), .IN2(search_data[21]), .S(
        \read_value_mux[12][21] ), .Q(n2245) );
  MUX21X1 U3413 ( .IN1(n1685), .IN2(search_data[8]), .S(
        \read_value_mux[12][8] ), .Q(n2244) );
  MUX21X1 U3414 ( .IN1(n1699), .IN2(search_data[13]), .S(
        \read_value_mux[12][13] ), .Q(n2243) );
  MUX21X1 U3415 ( .IN1(n1660), .IN2(search_data[0]), .S(
        \read_value_mux[12][0] ), .Q(n2242) );
  NAND4X0 U3416 ( .IN1(n2245), .IN2(n2244), .IN3(n2243), .IN4(n2242), .QN(
        n2246) );
  NOR4X0 U3417 ( .IN1(n2248), .IN2(n2247), .IN3(n1611), .IN4(n2246), .QN(n2270) );
  MUX21X1 U3418 ( .IN1(n1688), .IN2(search_data[9]), .S(
        \read_value_mux[12][9] ), .Q(n2252) );
  MUX21X1 U3419 ( .IN1(n1735), .IN2(search_data[29]), .S(
        \read_value_mux[12][29] ), .Q(n2251) );
  MUX21X1 U3420 ( .IN1(n1696), .IN2(search_data[12]), .S(
        \read_value_mux[12][12] ), .Q(n2250) );
  MUX21X1 U3421 ( .IN1(n1670), .IN2(search_data[3]), .S(
        \read_value_mux[12][3] ), .Q(n2249) );
  NAND4X0 U3422 ( .IN1(n2252), .IN2(n2251), .IN3(n2250), .IN4(n2249), .QN(
        n2268) );
  MUX21X1 U3423 ( .IN1(n1723), .IN2(search_data[22]), .S(
        \read_value_mux[12][22] ), .Q(n2256) );
  MUX21X1 U3424 ( .IN1(n1713), .IN2(search_data[18]), .S(
        \read_value_mux[12][18] ), .Q(n2255) );
  MUX21X1 U3425 ( .IN1(n1702), .IN2(search_data[14]), .S(
        \read_value_mux[12][14] ), .Q(n2254) );
  MUX21X1 U3426 ( .IN1(n1718), .IN2(search_data[20]), .S(
        \read_value_mux[12][20] ), .Q(n2253) );
  NAND4X0 U3427 ( .IN1(n2256), .IN2(n2255), .IN3(n2254), .IN4(n2253), .QN(
        n2267) );
  MUX21X1 U3428 ( .IN1(n1716), .IN2(search_data[19]), .S(
        \read_value_mux[12][19] ), .Q(n2260) );
  MUX21X1 U3429 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[12][24] ), .Q(n2259) );
  MUX21X1 U3430 ( .IN1(n1664), .IN2(search_data[1]), .S(
        \read_value_mux[12][1] ), .Q(n2258) );
  MUX21X1 U3431 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[12][23] ), .Q(n2257) );
  NAND4X0 U3432 ( .IN1(n2260), .IN2(n2259), .IN3(n2258), .IN4(n2257), .QN(
        n2266) );
  MUX21X1 U3433 ( .IN1(n1731), .IN2(search_data[27]), .S(
        \read_value_mux[12][27] ), .Q(n2264) );
  MUX21X1 U3434 ( .IN1(n1705), .IN2(n1704), .S(\read_value_mux[12][15] ), .Q(
        n2263) );
  MUX21X1 U3435 ( .IN1(n1673), .IN2(search_data[4]), .S(
        \read_value_mux[12][4] ), .Q(n2262) );
  MUX21X1 U3436 ( .IN1(n1740), .IN2(search_data[31]), .S(
        \read_value_mux[12][31] ), .Q(n2261) );
  NAND4X0 U3437 ( .IN1(n2264), .IN2(n2263), .IN3(n2262), .IN4(n2261), .QN(
        n2265) );
  NOR4X0 U3438 ( .IN1(n2268), .IN2(n2267), .IN3(n2266), .IN4(n2265), .QN(n2269) );
  NAND4X0 U3439 ( .IN1(n2272), .IN2(n2271), .IN3(n2270), .IN4(n2269), .QN(
        n3123) );
  NOR3X0 U3440 ( .IN1(n3064), .IN2(n3087), .IN3(n2923), .QN(n3008) );
  MUX21X1 U3441 ( .IN1(n1690), .IN2(n1691), .S(\read_value_mux[18][10] ), .Q(
        n2281) );
  MUX21X1 U3442 ( .IN1(search_data[4]), .IN2(n1672), .S(
        \read_value_mux[18][4] ), .Q(n2280) );
  MUX21X1 U3443 ( .IN1(search_data[21]), .IN2(n1719), .S(
        \read_value_mux[18][21] ), .Q(n2273) );
  AO221X1 U3444 ( .IN1(search_data[8]), .IN2(n1649), .IN3(n1686), .IN4(
        \read_value_mux[18][8] ), .IN5(n2273), .Q(n2279) );
  MUX21X1 U3445 ( .IN1(n1682), .IN2(search_data[7]), .S(
        \read_value_mux[18][7] ), .Q(n2276) );
  MUX21X1 U3446 ( .IN1(n1740), .IN2(search_data[31]), .S(
        \read_value_mux[18][31] ), .Q(n2275) );
  MUX21X1 U3447 ( .IN1(n1667), .IN2(search_data[2]), .S(
        \read_value_mux[18][2] ), .Q(n2274) );
  NAND4X0 U3448 ( .IN1(n2277), .IN2(n2276), .IN3(n2275), .IN4(n2274), .QN(
        n2278) );
  NOR4X0 U3449 ( .IN1(n2281), .IN2(n2280), .IN3(n2279), .IN4(n2278), .QN(n2313) );
  MUX21X1 U3450 ( .IN1(n1710), .IN2(search_data[17]), .S(
        \read_value_mux[18][17] ), .Q(n2282) );
  OA221X1 U3451 ( .IN1(search_data[27]), .IN2(n1652), .IN3(n1732), .IN4(
        \read_value_mux[18][27] ), .IN5(n2282), .Q(n2312) );
  MUX21X1 U3452 ( .IN1(search_data[30]), .IN2(n1737), .S(
        \read_value_mux[18][30] ), .Q(n2289) );
  MUX21X1 U3453 ( .IN1(search_data[13]), .IN2(n1698), .S(
        \read_value_mux[18][13] ), .Q(n2288) );
  MUX21X1 U3454 ( .IN1(n1718), .IN2(search_data[20]), .S(
        \read_value_mux[18][20] ), .Q(n2286) );
  MUX21X1 U3455 ( .IN1(n1735), .IN2(search_data[29]), .S(
        \read_value_mux[18][29] ), .Q(n2285) );
  MUX21X1 U3456 ( .IN1(n1670), .IN2(search_data[3]), .S(
        \read_value_mux[18][3] ), .Q(n2284) );
  MUX21X1 U3457 ( .IN1(n1729), .IN2(search_data[26]), .S(
        \read_value_mux[18][26] ), .Q(n2283) );
  NAND4X0 U3458 ( .IN1(n2286), .IN2(n2285), .IN3(n2284), .IN4(n2283), .QN(
        n2287) );
  NOR4X0 U3459 ( .IN1(n2289), .IN2(n2288), .IN3(n1611), .IN4(n2287), .QN(n2311) );
  MUX21X1 U3460 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[18][23] ), .Q(n2293) );
  MUX21X1 U3461 ( .IN1(n1707), .IN2(search_data[16]), .S(
        \read_value_mux[18][16] ), .Q(n2292) );
  MUX21X1 U3462 ( .IN1(n1679), .IN2(search_data[6]), .S(
        \read_value_mux[18][6] ), .Q(n2291) );
  MUX21X1 U3463 ( .IN1(n1688), .IN2(search_data[9]), .S(
        \read_value_mux[18][9] ), .Q(n2290) );
  NAND4X0 U3464 ( .IN1(n2293), .IN2(n2292), .IN3(n2291), .IN4(n2290), .QN(
        n2309) );
  MUX21X1 U3465 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[18][25] ), .Q(n2297) );
  MUX21X1 U3466 ( .IN1(n1723), .IN2(search_data[22]), .S(
        \read_value_mux[18][22] ), .Q(n2296) );
  MUX21X1 U3467 ( .IN1(n1694), .IN2(search_data[11]), .S(
        \read_value_mux[18][11] ), .Q(n2295) );
  MUX21X1 U3468 ( .IN1(n1714), .IN2(search_data[18]), .S(
        \read_value_mux[18][18] ), .Q(n2294) );
  NAND4X0 U3469 ( .IN1(n2297), .IN2(n2296), .IN3(n2295), .IN4(n2294), .QN(
        n2308) );
  MUX21X1 U3470 ( .IN1(n1716), .IN2(search_data[19]), .S(
        \read_value_mux[18][19] ), .Q(n2301) );
  MUX21X1 U3471 ( .IN1(n1660), .IN2(search_data[0]), .S(
        \read_value_mux[18][0] ), .Q(n2300) );
  MUX21X1 U3472 ( .IN1(n1676), .IN2(search_data[5]), .S(
        \read_value_mux[18][5] ), .Q(n2299) );
  MUX21X1 U3473 ( .IN1(n1702), .IN2(search_data[14]), .S(
        \read_value_mux[18][14] ), .Q(n2298) );
  NAND4X0 U3474 ( .IN1(n2301), .IN2(n2300), .IN3(n2299), .IN4(n2298), .QN(
        n2307) );
  MUX21X1 U3475 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[18][24] ), .Q(n2305) );
  MUX21X1 U3476 ( .IN1(n1696), .IN2(search_data[12]), .S(
        \read_value_mux[18][12] ), .Q(n2304) );
  MUX21X1 U3477 ( .IN1(n1664), .IN2(search_data[1]), .S(
        \read_value_mux[18][1] ), .Q(n2303) );
  MUX21X1 U3478 ( .IN1(n1705), .IN2(n1704), .S(\read_value_mux[18][15] ), .Q(
        n2302) );
  NAND4X0 U3479 ( .IN1(n2305), .IN2(n2304), .IN3(n2303), .IN4(n2302), .QN(
        n2306) );
  NOR4X0 U3480 ( .IN1(n2309), .IN2(n2308), .IN3(n2307), .IN4(n2306), .QN(n2310) );
  NAND4X0 U3481 ( .IN1(n2313), .IN2(n2312), .IN3(n2311), .IN4(n2310), .QN(
        n3082) );
  MUX21X1 U3482 ( .IN1(search_data[2]), .IN2(n1666), .S(
        \read_value_mux[20][2] ), .Q(n2322) );
  MUX21X1 U3483 ( .IN1(search_data[27]), .IN2(n1730), .S(
        \read_value_mux[20][27] ), .Q(n2321) );
  OAI22X1 U3484 ( .IN1(\read_value_mux[20][12] ), .IN2(n1697), .IN3(n1674), 
        .IN4(\read_value_mux[20][4] ), .QN(n2314) );
  AO221X1 U3485 ( .IN1(n1697), .IN2(\read_value_mux[20][12] ), .IN3(n1674), 
        .IN4(\read_value_mux[20][4] ), .IN5(n2314), .Q(n2320) );
  MUX21X1 U3486 ( .IN1(n1692), .IN2(n1690), .S(\read_value_mux[20][10] ), .Q(
        n2318) );
  MUX21X1 U3487 ( .IN1(n1723), .IN2(search_data[22]), .S(
        \read_value_mux[20][22] ), .Q(n2317) );
  MUX21X1 U3488 ( .IN1(n1707), .IN2(search_data[16]), .S(
        \read_value_mux[20][16] ), .Q(n2315) );
  NAND4X0 U3489 ( .IN1(n2318), .IN2(n2317), .IN3(n2316), .IN4(n2315), .QN(
        n2319) );
  NOR4X0 U3490 ( .IN1(n2322), .IN2(n2321), .IN3(n2320), .IN4(n2319), .QN(n2354) );
  AOI22X1 U3491 ( .IN1(n1741), .IN2(\read_value_mux[20][31] ), .IN3(n1727), 
        .IN4(\read_value_mux[20][25] ), .QN(n2323) );
  OA221X1 U3492 ( .IN1(n1741), .IN2(\read_value_mux[20][31] ), .IN3(n1727), 
        .IN4(\read_value_mux[20][25] ), .IN5(n2323), .Q(n2353) );
  MUX21X1 U3493 ( .IN1(search_data[17]), .IN2(n1709), .S(
        \read_value_mux[20][17] ), .Q(n2330) );
  MUX21X1 U3494 ( .IN1(search_data[8]), .IN2(n1684), .S(
        \read_value_mux[20][8] ), .Q(n2329) );
  MUX21X1 U3495 ( .IN1(n1699), .IN2(search_data[13]), .S(
        \read_value_mux[20][13] ), .Q(n2327) );
  MUX21X1 U3496 ( .IN1(n1682), .IN2(search_data[7]), .S(
        \read_value_mux[20][7] ), .Q(n2326) );
  MUX21X1 U3497 ( .IN1(n1712), .IN2(search_data[18]), .S(
        \read_value_mux[20][18] ), .Q(n2325) );
  MUX21X1 U3498 ( .IN1(n1688), .IN2(search_data[9]), .S(
        \read_value_mux[20][9] ), .Q(n2324) );
  NAND4X0 U3499 ( .IN1(n2327), .IN2(n2326), .IN3(n2325), .IN4(n2324), .QN(
        n2328) );
  NOR4X0 U3500 ( .IN1(n2330), .IN2(n2329), .IN3(n1611), .IN4(n2328), .QN(n2352) );
  MUX21X1 U3501 ( .IN1(n1705), .IN2(n1704), .S(\read_value_mux[20][15] ), .Q(
        n2334) );
  MUX21X1 U3502 ( .IN1(n1738), .IN2(search_data[30]), .S(
        \read_value_mux[20][30] ), .Q(n2333) );
  MUX21X1 U3503 ( .IN1(n1670), .IN2(search_data[3]), .S(
        \read_value_mux[20][3] ), .Q(n2332) );
  MUX21X1 U3504 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[20][24] ), .Q(n2331) );
  NAND4X0 U3505 ( .IN1(n2334), .IN2(n2333), .IN3(n2332), .IN4(n2331), .QN(
        n2350) );
  MUX21X1 U3506 ( .IN1(n1694), .IN2(search_data[11]), .S(
        \read_value_mux[20][11] ), .Q(n2338) );
  MUX21X1 U3507 ( .IN1(n1660), .IN2(search_data[0]), .S(
        \read_value_mux[20][0] ), .Q(n2337) );
  MUX21X1 U3508 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[20][23] ), .Q(n2336) );
  MUX21X1 U3509 ( .IN1(n1676), .IN2(search_data[5]), .S(
        \read_value_mux[20][5] ), .Q(n2335) );
  NAND4X0 U3510 ( .IN1(n2338), .IN2(n2337), .IN3(n2336), .IN4(n2335), .QN(
        n2349) );
  MUX21X1 U3511 ( .IN1(n1664), .IN2(search_data[1]), .S(
        \read_value_mux[20][1] ), .Q(n2342) );
  MUX21X1 U3512 ( .IN1(n1735), .IN2(search_data[29]), .S(
        \read_value_mux[20][29] ), .Q(n2341) );
  MUX21X1 U3513 ( .IN1(n1729), .IN2(search_data[26]), .S(
        \read_value_mux[20][26] ), .Q(n2340) );
  MUX21X1 U3514 ( .IN1(n1720), .IN2(search_data[21]), .S(
        \read_value_mux[20][21] ), .Q(n2339) );
  NAND4X0 U3515 ( .IN1(n2342), .IN2(n2341), .IN3(n2340), .IN4(n2339), .QN(
        n2348) );
  MUX21X1 U3516 ( .IN1(n1716), .IN2(search_data[19]), .S(
        \read_value_mux[20][19] ), .Q(n2346) );
  MUX21X1 U3517 ( .IN1(n1702), .IN2(search_data[14]), .S(
        \read_value_mux[20][14] ), .Q(n2345) );
  MUX21X1 U3518 ( .IN1(n1718), .IN2(search_data[20]), .S(
        \read_value_mux[20][20] ), .Q(n2344) );
  MUX21X1 U3519 ( .IN1(n1679), .IN2(search_data[6]), .S(
        \read_value_mux[20][6] ), .Q(n2343) );
  NAND4X0 U3520 ( .IN1(n2346), .IN2(n2345), .IN3(n2344), .IN4(n2343), .QN(
        n2347) );
  NOR4X0 U3521 ( .IN1(n2350), .IN2(n2349), .IN3(n2348), .IN4(n2347), .QN(n2351) );
  NAND4X0 U3522 ( .IN1(n2354), .IN2(n2353), .IN3(n2352), .IN4(n2351), .QN(
        n3067) );
  MUX21X1 U3523 ( .IN1(search_data[7]), .IN2(n1681), .S(
        \read_value_mux[21][7] ), .Q(n2395) );
  MUX21X1 U3524 ( .IN1(search_data[20]), .IN2(n1718), .S(
        \read_value_mux[21][20] ), .Q(n2394) );
  AOI22X1 U3525 ( .IN1(n1741), .IN2(\read_value_mux[21][31] ), .IN3(n1697), 
        .IN4(\read_value_mux[21][12] ), .QN(n2355) );
  OA221X1 U3526 ( .IN1(n1741), .IN2(\read_value_mux[21][31] ), .IN3(n1697), 
        .IN4(\read_value_mux[21][12] ), .IN5(n2355), .Q(n2360) );
  AOI22X1 U3527 ( .IN1(n1691), .IN2(\read_value_mux[21][10] ), .IN3(n1727), 
        .IN4(\read_value_mux[21][25] ), .QN(n2356) );
  OA221X1 U3528 ( .IN1(n1691), .IN2(\read_value_mux[21][10] ), .IN3(n1727), 
        .IN4(\read_value_mux[21][25] ), .IN5(n2356), .Q(n2359) );
  MUX21X1 U3529 ( .IN1(n1716), .IN2(search_data[19]), .S(
        \read_value_mux[21][19] ), .Q(n2358) );
  MUX21X1 U3530 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[21][24] ), .Q(n2357) );
  NAND4X0 U3531 ( .IN1(n2360), .IN2(n2359), .IN3(n2358), .IN4(n2357), .QN(
        n2393) );
  MUX21X1 U3532 ( .IN1(search_data[0]), .IN2(n1660), .S(
        \read_value_mux[21][0] ), .Q(n2367) );
  MUX21X1 U3533 ( .IN1(search_data[16]), .IN2(n1708), .S(
        \read_value_mux[21][16] ), .Q(n2366) );
  MUX21X1 U3534 ( .IN1(n1679), .IN2(search_data[6]), .S(
        \read_value_mux[21][6] ), .Q(n2364) );
  MUX21X1 U3535 ( .IN1(n1738), .IN2(search_data[30]), .S(
        \read_value_mux[21][30] ), .Q(n2363) );
  MUX21X1 U3536 ( .IN1(n1675), .IN2(search_data[5]), .S(
        \read_value_mux[21][5] ), .Q(n2362) );
  MUX21X1 U3537 ( .IN1(n1729), .IN2(search_data[26]), .S(
        \read_value_mux[21][26] ), .Q(n2361) );
  NAND4X0 U3538 ( .IN1(n2364), .IN2(n2363), .IN3(n2362), .IN4(n2361), .QN(
        n2365) );
  NOR4X0 U3539 ( .IN1(n2367), .IN2(n2366), .IN3(n1611), .IN4(n2365), .QN(n2391) );
  MUX21X1 U3540 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[21][23] ), .Q(n2371) );
  MUX21X1 U3541 ( .IN1(n1664), .IN2(search_data[1]), .S(
        \read_value_mux[21][1] ), .Q(n2370) );
  MUX21X1 U3542 ( .IN1(n1713), .IN2(search_data[18]), .S(
        \read_value_mux[21][18] ), .Q(n2369) );
  NAND4X0 U3543 ( .IN1(n2371), .IN2(n2370), .IN3(n2369), .IN4(n2368), .QN(
        n2387) );
  MUX21X1 U3544 ( .IN1(n1685), .IN2(search_data[8]), .S(
        \read_value_mux[21][8] ), .Q(n2375) );
  MUX21X1 U3545 ( .IN1(n1710), .IN2(search_data[17]), .S(
        \read_value_mux[21][17] ), .Q(n2374) );
  MUX21X1 U3546 ( .IN1(n1720), .IN2(search_data[21]), .S(
        \read_value_mux[21][21] ), .Q(n2373) );
  MUX21X1 U3547 ( .IN1(n1688), .IN2(search_data[9]), .S(
        \read_value_mux[21][9] ), .Q(n2372) );
  NAND4X0 U3548 ( .IN1(n2375), .IN2(n2374), .IN3(n2373), .IN4(n2372), .QN(
        n2386) );
  MUX21X1 U3549 ( .IN1(n1699), .IN2(search_data[13]), .S(
        \read_value_mux[21][13] ), .Q(n2379) );
  MUX21X1 U3550 ( .IN1(n1673), .IN2(search_data[4]), .S(
        \read_value_mux[21][4] ), .Q(n2378) );
  MUX21X1 U3551 ( .IN1(n1694), .IN2(search_data[11]), .S(
        \read_value_mux[21][11] ), .Q(n2377) );
  MUX21X1 U3552 ( .IN1(n1723), .IN2(search_data[22]), .S(
        \read_value_mux[21][22] ), .Q(n2376) );
  NAND4X0 U3553 ( .IN1(n2379), .IN2(n2378), .IN3(n2377), .IN4(n2376), .QN(
        n2385) );
  MUX21X1 U3554 ( .IN1(n1735), .IN2(search_data[29]), .S(
        \read_value_mux[21][29] ), .Q(n2383) );
  MUX21X1 U3555 ( .IN1(n1705), .IN2(n1704), .S(\read_value_mux[21][15] ), .Q(
        n2382) );
  MUX21X1 U3556 ( .IN1(n1667), .IN2(search_data[2]), .S(
        \read_value_mux[21][2] ), .Q(n2381) );
  MUX21X1 U3557 ( .IN1(n1702), .IN2(search_data[14]), .S(
        \read_value_mux[21][14] ), .Q(n2380) );
  NAND4X0 U3558 ( .IN1(n2383), .IN2(n2382), .IN3(n2381), .IN4(n2380), .QN(
        n2384) );
  NOR4X0 U3559 ( .IN1(n2387), .IN2(n2386), .IN3(n2385), .IN4(n2384), .QN(n2390) );
  MUX21X1 U3560 ( .IN1(n1731), .IN2(search_data[27]), .S(
        \read_value_mux[21][27] ), .Q(n2389) );
  MUX21X1 U3561 ( .IN1(n1670), .IN2(search_data[3]), .S(
        \read_value_mux[21][3] ), .Q(n2388) );
  NAND4X0 U3562 ( .IN1(n2391), .IN2(n2390), .IN3(n2389), .IN4(n2388), .QN(
        n2392) );
  NOR4X0 U3563 ( .IN1(n2395), .IN2(n2394), .IN3(n2393), .IN4(n2392), .QN(n3065) );
  MUX21X1 U3564 ( .IN1(search_data[13]), .IN2(n1698), .S(
        \read_value_mux[23][13] ), .Q(n2436) );
  MUX21X1 U3565 ( .IN1(search_data[7]), .IN2(n1681), .S(
        \read_value_mux[23][7] ), .Q(n2435) );
  AOI22X1 U3566 ( .IN1(n1695), .IN2(\read_value_mux[23][11] ), .IN3(n1708), 
        .IN4(\read_value_mux[23][16] ), .QN(n2396) );
  OA221X1 U3567 ( .IN1(n1695), .IN2(\read_value_mux[23][11] ), .IN3(n1708), 
        .IN4(\read_value_mux[23][16] ), .IN5(n2396), .Q(n2401) );
  AOI22X1 U3568 ( .IN1(n1725), .IN2(\read_value_mux[23][23] ), .IN3(n1671), 
        .IN4(\read_value_mux[23][3] ), .QN(n2397) );
  OA221X1 U3569 ( .IN1(n1725), .IN2(\read_value_mux[23][23] ), .IN3(n1671), 
        .IN4(\read_value_mux[23][3] ), .IN5(n2397), .Q(n2400) );
  MUX21X1 U3570 ( .IN1(n1692), .IN2(n1690), .S(\read_value_mux[23][10] ), .Q(
        n2399) );
  MUX21X1 U3571 ( .IN1(n1673), .IN2(search_data[4]), .S(
        \read_value_mux[23][4] ), .Q(n2398) );
  NAND4X0 U3572 ( .IN1(n2401), .IN2(n2400), .IN3(n2399), .IN4(n2398), .QN(
        n2434) );
  MUX21X1 U3573 ( .IN1(search_data[5]), .IN2(n1675), .S(
        \read_value_mux[23][5] ), .Q(n2408) );
  MUX21X1 U3574 ( .IN1(search_data[20]), .IN2(n1718), .S(
        \read_value_mux[23][20] ), .Q(n2407) );
  MUX21X1 U3575 ( .IN1(n1716), .IN2(search_data[19]), .S(
        \read_value_mux[23][19] ), .Q(n2405) );
  MUX21X1 U3576 ( .IN1(n1735), .IN2(search_data[29]), .S(
        \read_value_mux[23][29] ), .Q(n2404) );
  MUX21X1 U3577 ( .IN1(n1731), .IN2(search_data[27]), .S(
        \read_value_mux[23][27] ), .Q(n2403) );
  NAND4X0 U3578 ( .IN1(n2405), .IN2(n2404), .IN3(n2403), .IN4(n2402), .QN(
        n2406) );
  NOR4X0 U3579 ( .IN1(n2408), .IN2(n2407), .IN3(n1611), .IN4(n2406), .QN(n2432) );
  MUX21X1 U3580 ( .IN1(n1720), .IN2(search_data[21]), .S(
        \read_value_mux[23][21] ), .Q(n2412) );
  MUX21X1 U3581 ( .IN1(n1738), .IN2(search_data[30]), .S(
        \read_value_mux[23][30] ), .Q(n2411) );
  MUX21X1 U3582 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[23][25] ), .Q(n2410) );
  MUX21X1 U3583 ( .IN1(n1713), .IN2(search_data[18]), .S(
        \read_value_mux[23][18] ), .Q(n2409) );
  NAND4X0 U3584 ( .IN1(n2412), .IN2(n2411), .IN3(n2410), .IN4(n2409), .QN(
        n2428) );
  MUX21X1 U3585 ( .IN1(n1667), .IN2(search_data[2]), .S(
        \read_value_mux[23][2] ), .Q(n2416) );
  MUX21X1 U3586 ( .IN1(n1688), .IN2(search_data[9]), .S(
        \read_value_mux[23][9] ), .Q(n2415) );
  MUX21X1 U3587 ( .IN1(n1740), .IN2(search_data[31]), .S(
        \read_value_mux[23][31] ), .Q(n2414) );
  MUX21X1 U3588 ( .IN1(n1696), .IN2(search_data[12]), .S(
        \read_value_mux[23][12] ), .Q(n2413) );
  NAND4X0 U3589 ( .IN1(n2416), .IN2(n2415), .IN3(n2414), .IN4(n2413), .QN(
        n2427) );
  MUX21X1 U3590 ( .IN1(n1661), .IN2(search_data[0]), .S(
        \read_value_mux[23][0] ), .Q(n2420) );
  MUX21X1 U3591 ( .IN1(n1729), .IN2(search_data[26]), .S(
        \read_value_mux[23][26] ), .Q(n2419) );
  MUX21X1 U3592 ( .IN1(n1723), .IN2(search_data[22]), .S(
        \read_value_mux[23][22] ), .Q(n2418) );
  MUX21X1 U3593 ( .IN1(n1702), .IN2(search_data[14]), .S(
        \read_value_mux[23][14] ), .Q(n2417) );
  NAND4X0 U3594 ( .IN1(n2420), .IN2(n2419), .IN3(n2418), .IN4(n2417), .QN(
        n2426) );
  MUX21X1 U3595 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[23][24] ), .Q(n2424) );
  MUX21X1 U3596 ( .IN1(n1710), .IN2(search_data[17]), .S(
        \read_value_mux[23][17] ), .Q(n2423) );
  MUX21X1 U3597 ( .IN1(n1684), .IN2(search_data[8]), .S(
        \read_value_mux[23][8] ), .Q(n2422) );
  MUX21X1 U3598 ( .IN1(n1679), .IN2(search_data[6]), .S(
        \read_value_mux[23][6] ), .Q(n2421) );
  NAND4X0 U3599 ( .IN1(n2424), .IN2(n2423), .IN3(n2422), .IN4(n2421), .QN(
        n2425) );
  NOR4X0 U3600 ( .IN1(n2428), .IN2(n2427), .IN3(n2426), .IN4(n2425), .QN(n2431) );
  MUX21X1 U3601 ( .IN1(n1705), .IN2(n1704), .S(\read_value_mux[23][15] ), .Q(
        n2430) );
  MUX21X1 U3602 ( .IN1(n1664), .IN2(search_data[1]), .S(
        \read_value_mux[23][1] ), .Q(n2429) );
  NAND4X0 U3603 ( .IN1(n2432), .IN2(n2431), .IN3(n2430), .IN4(n2429), .QN(
        n2433) );
  NOR4X0 U3604 ( .IN1(n2436), .IN2(n2435), .IN3(n2434), .IN4(n2433), .QN(n3068) );
  MUX21X1 U3605 ( .IN1(search_data[7]), .IN2(n1681), .S(
        \read_value_mux[24][7] ), .Q(n2445) );
  MUX21X1 U3606 ( .IN1(search_data[21]), .IN2(n1719), .S(
        \read_value_mux[24][21] ), .Q(n2444) );
  OAI22X1 U3607 ( .IN1(n1711), .IN2(\read_value_mux[24][17] ), .IN3(n1661), 
        .IN4(\read_value_mux[24][0] ), .QN(n2437) );
  AO221X1 U3608 ( .IN1(n1711), .IN2(\read_value_mux[24][17] ), .IN3(
        \read_value_mux[24][0] ), .IN4(n1661), .IN5(n2437), .Q(n2443) );
  MUX21X1 U3609 ( .IN1(n1735), .IN2(search_data[29]), .S(
        \read_value_mux[24][29] ), .Q(n2441) );
  MUX21X1 U3610 ( .IN1(n1707), .IN2(search_data[16]), .S(
        \read_value_mux[24][16] ), .Q(n2440) );
  MUX21X1 U3611 ( .IN1(n1679), .IN2(search_data[6]), .S(
        \read_value_mux[24][6] ), .Q(n2439) );
  MUX21X1 U3612 ( .IN1(n1670), .IN2(search_data[3]), .S(
        \read_value_mux[24][3] ), .Q(n2438) );
  NAND4X0 U3613 ( .IN1(n2441), .IN2(n2440), .IN3(n2439), .IN4(n2438), .QN(
        n2442) );
  NOR4X0 U3614 ( .IN1(n2445), .IN2(n2444), .IN3(n2443), .IN4(n2442), .QN(n2477) );
  AOI22X1 U3615 ( .IN1(n1703), .IN2(\read_value_mux[24][14] ), .IN3(n1739), 
        .IN4(\read_value_mux[24][30] ), .QN(n2446) );
  OA221X1 U3616 ( .IN1(n1703), .IN2(\read_value_mux[24][14] ), .IN3(n1739), 
        .IN4(\read_value_mux[24][30] ), .IN5(n2446), .Q(n2476) );
  MUX21X1 U3617 ( .IN1(n1704), .IN2(n1705), .S(\read_value_mux[24][15] ), .Q(
        n2453) );
  MUX21X1 U3618 ( .IN1(search_data[13]), .IN2(n1698), .S(
        \read_value_mux[24][13] ), .Q(n2452) );
  MUX21X1 U3619 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[24][23] ), .Q(n2450) );
  MUX21X1 U3620 ( .IN1(n1692), .IN2(n1690), .S(\read_value_mux[24][10] ), .Q(
        n2449) );
  MUX21X1 U3621 ( .IN1(n1723), .IN2(search_data[22]), .S(
        \read_value_mux[24][22] ), .Q(n2448) );
  MUX21X1 U3622 ( .IN1(n1729), .IN2(search_data[26]), .S(
        \read_value_mux[24][26] ), .Q(n2447) );
  NAND4X0 U3623 ( .IN1(n2450), .IN2(n2449), .IN3(n2448), .IN4(n2447), .QN(
        n2451) );
  NOR4X0 U3624 ( .IN1(n2453), .IN2(n2452), .IN3(n1611), .IN4(n2451), .QN(n2475) );
  MUX21X1 U3625 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[24][28] ), .Q(n2457) );
  MUX21X1 U3626 ( .IN1(n1667), .IN2(search_data[2]), .S(
        \read_value_mux[24][2] ), .Q(n2456) );
  MUX21X1 U3627 ( .IN1(n1673), .IN2(search_data[4]), .S(
        \read_value_mux[24][4] ), .Q(n2455) );
  MUX21X1 U3628 ( .IN1(n1741), .IN2(search_data[31]), .S(
        \read_value_mux[24][31] ), .Q(n2454) );
  NAND4X0 U3629 ( .IN1(n2457), .IN2(n2456), .IN3(n2455), .IN4(n2454), .QN(
        n2473) );
  MUX21X1 U3630 ( .IN1(n1684), .IN2(search_data[8]), .S(
        \read_value_mux[24][8] ), .Q(n2461) );
  MUX21X1 U3631 ( .IN1(n1716), .IN2(search_data[19]), .S(
        \read_value_mux[24][19] ), .Q(n2460) );
  MUX21X1 U3632 ( .IN1(n1688), .IN2(search_data[9]), .S(
        \read_value_mux[24][9] ), .Q(n2459) );
  MUX21X1 U3633 ( .IN1(n1713), .IN2(search_data[18]), .S(
        \read_value_mux[24][18] ), .Q(n2458) );
  NAND4X0 U3634 ( .IN1(n2461), .IN2(n2460), .IN3(n2459), .IN4(n2458), .QN(
        n2472) );
  MUX21X1 U3635 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[24][25] ), .Q(n2465) );
  MUX21X1 U3636 ( .IN1(n1718), .IN2(search_data[20]), .S(
        \read_value_mux[24][20] ), .Q(n2464) );
  MUX21X1 U3637 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[24][24] ), .Q(n2463) );
  MUX21X1 U3638 ( .IN1(n1694), .IN2(search_data[11]), .S(
        \read_value_mux[24][11] ), .Q(n2462) );
  NAND4X0 U3639 ( .IN1(n2465), .IN2(n2464), .IN3(n2463), .IN4(n2462), .QN(
        n2471) );
  MUX21X1 U3640 ( .IN1(n1664), .IN2(search_data[1]), .S(
        \read_value_mux[24][1] ), .Q(n2469) );
  MUX21X1 U3641 ( .IN1(n1731), .IN2(search_data[27]), .S(
        \read_value_mux[24][27] ), .Q(n2468) );
  MUX21X1 U3642 ( .IN1(n1675), .IN2(search_data[5]), .S(
        \read_value_mux[24][5] ), .Q(n2467) );
  MUX21X1 U3643 ( .IN1(n1696), .IN2(search_data[12]), .S(
        \read_value_mux[24][12] ), .Q(n2466) );
  NAND4X0 U3644 ( .IN1(n2469), .IN2(n2468), .IN3(n2467), .IN4(n2466), .QN(
        n2470) );
  NOR4X0 U3645 ( .IN1(n2473), .IN2(n2472), .IN3(n2471), .IN4(n2470), .QN(n2474) );
  NAND4X0 U3646 ( .IN1(n2477), .IN2(n2476), .IN3(n2475), .IN4(n2474), .QN(
        n3111) );
  MUX21X1 U3647 ( .IN1(search_data[16]), .IN2(n1708), .S(
        \read_value_mux[26][16] ), .Q(n2486) );
  MUX21X1 U3648 ( .IN1(search_data[24]), .IN2(n1726), .S(
        \read_value_mux[26][24] ), .Q(n2485) );
  OAI22X1 U3649 ( .IN1(\read_value_mux[26][17] ), .IN2(n1711), .IN3(n1695), 
        .IN4(\read_value_mux[26][11] ), .QN(n2478) );
  AO221X1 U3650 ( .IN1(n1711), .IN2(\read_value_mux[26][17] ), .IN3(n1695), 
        .IN4(\read_value_mux[26][11] ), .IN5(n2478), .Q(n2484) );
  MUX21X1 U3651 ( .IN1(n1699), .IN2(search_data[13]), .S(
        \read_value_mux[26][13] ), .Q(n2482) );
  MUX21X1 U3652 ( .IN1(n1705), .IN2(n1704), .S(\read_value_mux[26][15] ), .Q(
        n2481) );
  MUX21X1 U3653 ( .IN1(n1684), .IN2(search_data[8]), .S(
        \read_value_mux[26][8] ), .Q(n2480) );
  MUX21X1 U3654 ( .IN1(n1692), .IN2(search_data[10]), .S(
        \read_value_mux[26][10] ), .Q(n2479) );
  NAND4X0 U3655 ( .IN1(n2482), .IN2(n2481), .IN3(n2480), .IN4(n2479), .QN(
        n2483) );
  NOR4X0 U3656 ( .IN1(n2486), .IN2(n2485), .IN3(n2484), .IN4(n2483), .QN(n2518) );
  MUX21X1 U3657 ( .IN1(n1696), .IN2(search_data[12]), .S(
        \read_value_mux[26][12] ), .Q(n2487) );
  OA221X1 U3658 ( .IN1(search_data[21]), .IN2(n1653), .IN3(n1721), .IN4(
        \read_value_mux[26][21] ), .IN5(n2487), .Q(n2517) );
  MUX21X1 U3659 ( .IN1(search_data[3]), .IN2(n1669), .S(
        \read_value_mux[26][3] ), .Q(n2494) );
  MUX21X1 U3660 ( .IN1(search_data[9]), .IN2(n1687), .S(
        \read_value_mux[26][9] ), .Q(n2493) );
  MUX21X1 U3661 ( .IN1(n1682), .IN2(search_data[7]), .S(
        \read_value_mux[26][7] ), .Q(n2491) );
  MUX21X1 U3662 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[26][28] ), .Q(n2490) );
  MUX21X1 U3663 ( .IN1(n1731), .IN2(search_data[27]), .S(
        \read_value_mux[26][27] ), .Q(n2489) );
  MUX21X1 U3664 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[26][25] ), .Q(n2488) );
  NAND4X0 U3665 ( .IN1(n2491), .IN2(n2490), .IN3(n2489), .IN4(n2488), .QN(
        n2492) );
  NOR4X0 U3666 ( .IN1(n2494), .IN2(n2493), .IN3(n1611), .IN4(n2492), .QN(n2516) );
  MUX21X1 U3667 ( .IN1(n1702), .IN2(search_data[14]), .S(
        \read_value_mux[26][14] ), .Q(n2498) );
  MUX21X1 U3668 ( .IN1(n1716), .IN2(search_data[19]), .S(
        \read_value_mux[26][19] ), .Q(n2497) );
  MUX21X1 U3669 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[26][23] ), .Q(n2496) );
  MUX21X1 U3670 ( .IN1(n1718), .IN2(search_data[20]), .S(
        \read_value_mux[26][20] ), .Q(n2495) );
  NAND4X0 U3671 ( .IN1(n2498), .IN2(n2497), .IN3(n2496), .IN4(n2495), .QN(
        n2514) );
  MUX21X1 U3672 ( .IN1(n1723), .IN2(search_data[22]), .S(
        \read_value_mux[26][22] ), .Q(n2502) );
  MUX21X1 U3673 ( .IN1(n1664), .IN2(search_data[1]), .S(
        \read_value_mux[26][1] ), .Q(n2501) );
  MUX21X1 U3674 ( .IN1(n1679), .IN2(search_data[6]), .S(
        \read_value_mux[26][6] ), .Q(n2500) );
  MUX21X1 U3675 ( .IN1(n1673), .IN2(search_data[4]), .S(
        \read_value_mux[26][4] ), .Q(n2499) );
  NAND4X0 U3676 ( .IN1(n2502), .IN2(n2501), .IN3(n2500), .IN4(n2499), .QN(
        n2513) );
  MUX21X1 U3677 ( .IN1(n1738), .IN2(search_data[30]), .S(
        \read_value_mux[26][30] ), .Q(n2506) );
  MUX21X1 U3678 ( .IN1(n1735), .IN2(search_data[29]), .S(
        \read_value_mux[26][29] ), .Q(n2505) );
  MUX21X1 U3679 ( .IN1(n1675), .IN2(search_data[5]), .S(
        \read_value_mux[26][5] ), .Q(n2504) );
  MUX21X1 U3680 ( .IN1(n1729), .IN2(search_data[26]), .S(
        \read_value_mux[26][26] ), .Q(n2503) );
  NAND4X0 U3681 ( .IN1(n2506), .IN2(n2505), .IN3(n2504), .IN4(n2503), .QN(
        n2512) );
  MUX21X1 U3682 ( .IN1(n1667), .IN2(search_data[2]), .S(
        \read_value_mux[26][2] ), .Q(n2510) );
  MUX21X1 U3683 ( .IN1(n1740), .IN2(search_data[31]), .S(
        \read_value_mux[26][31] ), .Q(n2509) );
  MUX21X1 U3684 ( .IN1(n1661), .IN2(search_data[0]), .S(
        \read_value_mux[26][0] ), .Q(n2508) );
  MUX21X1 U3685 ( .IN1(n1713), .IN2(search_data[18]), .S(
        \read_value_mux[26][18] ), .Q(n2507) );
  NAND4X0 U3686 ( .IN1(n2510), .IN2(n2509), .IN3(n2508), .IN4(n2507), .QN(
        n2511) );
  NOR4X0 U3687 ( .IN1(n2514), .IN2(n2513), .IN3(n2512), .IN4(n2511), .QN(n2515) );
  NAND4X0 U3688 ( .IN1(n2518), .IN2(n2517), .IN3(n2516), .IN4(n2515), .QN(
        n3071) );
  OAI22X1 U3689 ( .IN1(\read_value_mux[27][5] ), .IN2(n1677), .IN3(n1689), 
        .IN4(\read_value_mux[27][9] ), .QN(n2519) );
  AO221X1 U3690 ( .IN1(n1677), .IN2(\read_value_mux[27][5] ), .IN3(n1689), 
        .IN4(\read_value_mux[27][9] ), .IN5(n2519), .Q(n2559) );
  OAI22X1 U3691 ( .IN1(\read_value_mux[27][18] ), .IN2(n1713), .IN3(n1741), 
        .IN4(\read_value_mux[27][31] ), .QN(n2520) );
  AO221X1 U3692 ( .IN1(n1712), .IN2(\read_value_mux[27][18] ), .IN3(n1741), 
        .IN4(\read_value_mux[27][31] ), .IN5(n2520), .Q(n2558) );
  MUX21X1 U3693 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[27][23] ), .Q(n2524) );
  MUX21X1 U3694 ( .IN1(n1699), .IN2(search_data[13]), .S(
        \read_value_mux[27][13] ), .Q(n2523) );
  MUX21X1 U3695 ( .IN1(n1697), .IN2(search_data[12]), .S(
        \read_value_mux[27][12] ), .Q(n2522) );
  MUX21X1 U3696 ( .IN1(n1692), .IN2(search_data[10]), .S(
        \read_value_mux[27][10] ), .Q(n2521) );
  NAND4X0 U3697 ( .IN1(n2524), .IN2(n2523), .IN3(n2522), .IN4(n2521), .QN(
        n2557) );
  MUX21X1 U3698 ( .IN1(search_data[14]), .IN2(n1701), .S(
        \read_value_mux[27][14] ), .Q(n2531) );
  MUX21X1 U3699 ( .IN1(search_data[19]), .IN2(n1716), .S(
        \read_value_mux[27][19] ), .Q(n2530) );
  MUX21X1 U3700 ( .IN1(n1731), .IN2(search_data[27]), .S(
        \read_value_mux[27][27] ), .Q(n2528) );
  MUX21X1 U3701 ( .IN1(n1682), .IN2(search_data[7]), .S(
        \read_value_mux[27][7] ), .Q(n2527) );
  MUX21X1 U3702 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[27][25] ), .Q(n2526) );
  MUX21X1 U3703 ( .IN1(n1707), .IN2(search_data[16]), .S(
        \read_value_mux[27][16] ), .Q(n2525) );
  NAND4X0 U3704 ( .IN1(n2528), .IN2(n2527), .IN3(n2526), .IN4(n2525), .QN(
        n2529) );
  NOR4X0 U3705 ( .IN1(n2531), .IN2(n2530), .IN3(n1611), .IN4(n2529), .QN(n2555) );
  MUX21X1 U3706 ( .IN1(n1710), .IN2(search_data[17]), .S(
        \read_value_mux[27][17] ), .Q(n2535) );
  MUX21X1 U3707 ( .IN1(n1669), .IN2(search_data[3]), .S(
        \read_value_mux[27][3] ), .Q(n2534) );
  MUX21X1 U3708 ( .IN1(n1738), .IN2(search_data[30]), .S(
        \read_value_mux[27][30] ), .Q(n2533) );
  MUX21X1 U3709 ( .IN1(n1663), .IN2(search_data[1]), .S(
        \read_value_mux[27][1] ), .Q(n2532) );
  NAND4X0 U3710 ( .IN1(n2535), .IN2(n2534), .IN3(n2533), .IN4(n2532), .QN(
        n2551) );
  MUX21X1 U3711 ( .IN1(n1729), .IN2(search_data[26]), .S(
        \read_value_mux[27][26] ), .Q(n2539) );
  MUX21X1 U3712 ( .IN1(n1705), .IN2(n1704), .S(\read_value_mux[27][15] ), .Q(
        n2538) );
  MUX21X1 U3713 ( .IN1(n1694), .IN2(search_data[11]), .S(
        \read_value_mux[27][11] ), .Q(n2537) );
  MUX21X1 U3714 ( .IN1(n1660), .IN2(search_data[0]), .S(
        \read_value_mux[27][0] ), .Q(n2536) );
  NAND4X0 U3715 ( .IN1(n2539), .IN2(n2538), .IN3(n2537), .IN4(n2536), .QN(
        n2550) );
  MUX21X1 U3716 ( .IN1(n1722), .IN2(search_data[22]), .S(
        \read_value_mux[27][22] ), .Q(n2543) );
  MUX21X1 U3717 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[27][24] ), .Q(n2542) );
  MUX21X1 U3718 ( .IN1(n1679), .IN2(search_data[6]), .S(
        \read_value_mux[27][6] ), .Q(n2541) );
  MUX21X1 U3719 ( .IN1(n1735), .IN2(search_data[29]), .S(
        \read_value_mux[27][29] ), .Q(n2540) );
  NAND4X0 U3720 ( .IN1(n2543), .IN2(n2542), .IN3(n2541), .IN4(n2540), .QN(
        n2549) );
  MUX21X1 U3721 ( .IN1(n1718), .IN2(search_data[20]), .S(
        \read_value_mux[27][20] ), .Q(n2547) );
  MUX21X1 U3722 ( .IN1(n1684), .IN2(search_data[8]), .S(
        \read_value_mux[27][8] ), .Q(n2546) );
  MUX21X1 U3723 ( .IN1(n1666), .IN2(search_data[2]), .S(
        \read_value_mux[27][2] ), .Q(n2545) );
  MUX21X1 U3724 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[27][28] ), .Q(n2544) );
  NAND4X0 U3725 ( .IN1(n2547), .IN2(n2546), .IN3(n2545), .IN4(n2544), .QN(
        n2548) );
  NOR4X0 U3726 ( .IN1(n2551), .IN2(n2550), .IN3(n2549), .IN4(n2548), .QN(n2554) );
  MUX21X1 U3727 ( .IN1(n1673), .IN2(search_data[4]), .S(
        \read_value_mux[27][4] ), .Q(n2553) );
  MUX21X1 U3728 ( .IN1(n1720), .IN2(search_data[21]), .S(
        \read_value_mux[27][21] ), .Q(n2552) );
  NAND4X0 U3729 ( .IN1(n2554), .IN2(n2555), .IN3(n2553), .IN4(n2552), .QN(
        n2556) );
  NOR4X0 U3730 ( .IN1(n2556), .IN2(n2558), .IN3(n2557), .IN4(n2559), .QN(n3072) );
  MUX21X1 U3731 ( .IN1(search_data[19]), .IN2(n1716), .S(
        \read_value_mux[29][19] ), .Q(n2593) );
  MUX21X1 U3732 ( .IN1(search_data[31]), .IN2(n1740), .S(
        \read_value_mux[29][31] ), .Q(n2592) );
  AOI22X1 U3733 ( .IN1(n1732), .IN2(\read_value_mux[29][27] ), .IN3(n1736), 
        .IN4(\read_value_mux[29][29] ), .QN(n2560) );
  OA221X1 U3734 ( .IN1(n1732), .IN2(\read_value_mux[29][27] ), .IN3(n1736), 
        .IN4(\read_value_mux[29][29] ), .IN5(n2560), .Q(n2565) );
  AOI22X1 U3735 ( .IN1(n1677), .IN2(\read_value_mux[29][5] ), .IN3(n1718), 
        .IN4(\read_value_mux[29][20] ), .QN(n2561) );
  OA221X1 U3736 ( .IN1(n1677), .IN2(\read_value_mux[29][5] ), .IN3(n1718), 
        .IN4(\read_value_mux[29][20] ), .IN5(n2561), .Q(n2564) );
  MUX21X1 U3737 ( .IN1(n1705), .IN2(n1704), .S(\read_value_mux[29][15] ), .Q(
        n2563) );
  MUX21X1 U3738 ( .IN1(n1663), .IN2(search_data[1]), .S(
        \read_value_mux[29][1] ), .Q(n2562) );
  MUX21X1 U3739 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[29][28] ), .Q(n2567) );
  MUX21X1 U3740 ( .IN1(n1699), .IN2(search_data[13]), .S(
        \read_value_mux[29][13] ), .Q(n2566) );
  MUX21X1 U3741 ( .IN1(n1719), .IN2(search_data[21]), .S(
        \read_value_mux[29][21] ), .Q(n2571) );
  MUX21X1 U3742 ( .IN1(n1729), .IN2(search_data[26]), .S(
        \read_value_mux[29][26] ), .Q(n2570) );
  MUX21X1 U3743 ( .IN1(n1685), .IN2(search_data[8]), .S(
        \read_value_mux[29][8] ), .Q(n2569) );
  NAND4X0 U3744 ( .IN1(n2571), .IN2(n2570), .IN3(n2569), .IN4(n2568), .QN(
        n2587) );
  MUX21X1 U3745 ( .IN1(n1697), .IN2(search_data[12]), .S(
        \read_value_mux[29][12] ), .Q(n2574) );
  MUX21X1 U3746 ( .IN1(n1738), .IN2(search_data[30]), .S(
        \read_value_mux[29][30] ), .Q(n2573) );
  MUX21X1 U3747 ( .IN1(n1667), .IN2(search_data[2]), .S(
        \read_value_mux[29][2] ), .Q(n2572) );
  NAND4X0 U3748 ( .IN1(n2575), .IN2(n2574), .IN3(n2573), .IN4(n2572), .QN(
        n2586) );
  MUX21X1 U3749 ( .IN1(n1710), .IN2(search_data[17]), .S(
        \read_value_mux[29][17] ), .Q(n2579) );
  MUX21X1 U3750 ( .IN1(n1714), .IN2(search_data[18]), .S(
        \read_value_mux[29][18] ), .Q(n2578) );
  MUX21X1 U3751 ( .IN1(n1702), .IN2(search_data[14]), .S(
        \read_value_mux[29][14] ), .Q(n2576) );
  NAND4X0 U3752 ( .IN1(n2579), .IN2(n2578), .IN3(n2577), .IN4(n2576), .QN(
        n2585) );
  MUX21X1 U3753 ( .IN1(n1678), .IN2(search_data[6]), .S(
        \read_value_mux[29][6] ), .Q(n2583) );
  MUX21X1 U3754 ( .IN1(n1669), .IN2(search_data[3]), .S(
        \read_value_mux[29][3] ), .Q(n2581) );
  MUX21X1 U3755 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[29][25] ), .Q(n2580) );
  NAND4X0 U3756 ( .IN1(n2583), .IN2(n2582), .IN3(n2581), .IN4(n2580), .QN(
        n2584) );
  MUX21X1 U3757 ( .IN1(n1694), .IN2(search_data[11]), .S(
        \read_value_mux[29][11] ), .Q(n2589) );
  MUX21X1 U3758 ( .IN1(n1707), .IN2(search_data[16]), .S(
        \read_value_mux[29][16] ), .Q(n2588) );
  OAI22X1 U3759 ( .IN1(\read_value_mux[31][7] ), .IN2(n1683), .IN3(n1674), 
        .IN4(\read_value_mux[31][4] ), .QN(n2594) );
  MUX21X1 U3760 ( .IN1(n1702), .IN2(search_data[14]), .S(
        \read_value_mux[31][14] ), .Q(n2598) );
  MUX21X1 U3761 ( .IN1(n1666), .IN2(search_data[2]), .S(
        \read_value_mux[31][2] ), .Q(n2597) );
  MUX21X1 U3762 ( .IN1(n1731), .IN2(search_data[27]), .S(
        \read_value_mux[31][27] ), .Q(n2596) );
  MUX21X1 U3763 ( .IN1(n1696), .IN2(search_data[12]), .S(
        \read_value_mux[31][12] ), .Q(n2595) );
  NAND4X0 U3764 ( .IN1(n2598), .IN2(n2597), .IN3(n2596), .IN4(n2595), .QN(
        n2631) );
  MUX21X1 U3765 ( .IN1(search_data[24]), .IN2(n1726), .S(
        \read_value_mux[31][24] ), .Q(n2605) );
  MUX21X1 U3766 ( .IN1(search_data[17]), .IN2(n1709), .S(
        \read_value_mux[31][17] ), .Q(n2604) );
  MUX21X1 U3767 ( .IN1(n1678), .IN2(search_data[6]), .S(
        \read_value_mux[31][6] ), .Q(n2602) );
  MUX21X1 U3768 ( .IN1(n1741), .IN2(search_data[31]), .S(
        \read_value_mux[31][31] ), .Q(n2601) );
  MUX21X1 U3769 ( .IN1(n1722), .IN2(search_data[22]), .S(
        \read_value_mux[31][22] ), .Q(n2600) );
  NAND4X0 U3770 ( .IN1(n2602), .IN2(n2601), .IN3(n2600), .IN4(n2599), .QN(
        n2603) );
  MUX21X1 U3771 ( .IN1(n1735), .IN2(search_data[29]), .S(
        \read_value_mux[31][29] ), .Q(n2609) );
  MUX21X1 U3772 ( .IN1(n1662), .IN2(search_data[0]), .S(
        \read_value_mux[31][0] ), .Q(n2607) );
  MUX21X1 U3773 ( .IN1(n1712), .IN2(search_data[18]), .S(
        \read_value_mux[31][18] ), .Q(n2606) );
  NAND4X0 U3774 ( .IN1(n2609), .IN2(n2608), .IN3(n2607), .IN4(n2606), .QN(
        n2625) );
  MUX21X1 U3775 ( .IN1(n1663), .IN2(search_data[1]), .S(
        \read_value_mux[31][1] ), .Q(n2613) );
  MUX21X1 U3776 ( .IN1(n1688), .IN2(search_data[9]), .S(
        \read_value_mux[31][9] ), .Q(n2612) );
  MUX21X1 U3777 ( .IN1(n1698), .IN2(search_data[13]), .S(
        \read_value_mux[31][13] ), .Q(n2610) );
  NAND4X0 U3778 ( .IN1(n2613), .IN2(n2612), .IN3(n2611), .IN4(n2610), .QN(
        n2624) );
  MUX21X1 U3779 ( .IN1(n1715), .IN2(search_data[19]), .S(
        \read_value_mux[31][19] ), .Q(n2617) );
  MUX21X1 U3780 ( .IN1(n1706), .IN2(n1704), .S(\read_value_mux[31][15] ), .Q(
        n2616) );
  MUX21X1 U3781 ( .IN1(n1707), .IN2(search_data[16]), .S(
        \read_value_mux[31][16] ), .Q(n2614) );
  NAND4X0 U3782 ( .IN1(n2617), .IN2(n2616), .IN3(n2615), .IN4(n2614), .QN(
        n2623) );
  MUX21X1 U3783 ( .IN1(n1720), .IN2(search_data[21]), .S(
        \read_value_mux[31][21] ), .Q(n2621) );
  MUX21X1 U3784 ( .IN1(n1737), .IN2(search_data[30]), .S(
        \read_value_mux[31][30] ), .Q(n2618) );
  NAND4X0 U3785 ( .IN1(n2621), .IN2(n2620), .IN3(n2619), .IN4(n2618), .QN(
        n2622) );
  NOR4X0 U3786 ( .IN1(n2625), .IN2(n2624), .IN3(n2623), .IN4(n2622), .QN(n2628) );
  MUX21X1 U3787 ( .IN1(n1675), .IN2(search_data[5]), .S(
        \read_value_mux[31][5] ), .Q(n2627) );
  MUX21X1 U3788 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[31][28] ), .Q(n2626) );
  NAND4X0 U3789 ( .IN1(n2629), .IN2(n2628), .IN3(n2627), .IN4(n2626), .QN(
        n2630) );
  MUX21X1 U3790 ( .IN1(search_data[9]), .IN2(n1687), .S(
        \read_value_mux[30][9] ), .Q(n2642) );
  MUX21X1 U3791 ( .IN1(search_data[14]), .IN2(n1701), .S(
        \read_value_mux[30][14] ), .Q(n2641) );
  OAI22X1 U3792 ( .IN1(n1677), .IN2(\read_value_mux[30][5] ), .IN3(n1706), 
        .IN4(\read_value_mux[30][15] ), .QN(n2634) );
  AO221X1 U3793 ( .IN1(n1677), .IN2(\read_value_mux[30][5] ), .IN3(
        \read_value_mux[30][15] ), .IN4(n1706), .IN5(n2634), .Q(n2640) );
  MUX21X1 U3794 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[30][28] ), .Q(n2638) );
  MUX21X1 U3795 ( .IN1(n1681), .IN2(search_data[7]), .S(
        \read_value_mux[30][7] ), .Q(n2637) );
  MUX21X1 U3796 ( .IN1(n1684), .IN2(search_data[8]), .S(
        \read_value_mux[30][8] ), .Q(n2636) );
  MUX21X1 U3797 ( .IN1(n1740), .IN2(search_data[31]), .S(
        \read_value_mux[30][31] ), .Q(n2635) );
  NAND4X0 U3798 ( .IN1(n2638), .IN2(n2637), .IN3(n2636), .IN4(n2635), .QN(
        n2639) );
  NOR4X0 U3799 ( .IN1(n2642), .IN2(n2641), .IN3(n2640), .IN4(n2639), .QN(n2674) );
  AOI22X1 U3800 ( .IN1(n1668), .IN2(\read_value_mux[30][2] ), .IN3(n1671), 
        .IN4(\read_value_mux[30][3] ), .QN(n2643) );
  OA221X1 U3801 ( .IN1(n1668), .IN2(\read_value_mux[30][2] ), .IN3(n1671), 
        .IN4(\read_value_mux[30][3] ), .IN5(n2643), .Q(n2673) );
  MUX21X1 U3802 ( .IN1(search_data[22]), .IN2(n1722), .S(
        \read_value_mux[30][22] ), .Q(n2650) );
  MUX21X1 U3803 ( .IN1(search_data[24]), .IN2(n1726), .S(
        \read_value_mux[30][24] ), .Q(n2649) );
  MUX21X1 U3804 ( .IN1(n1728), .IN2(search_data[26]), .S(
        \read_value_mux[30][26] ), .Q(n2647) );
  MUX21X1 U3805 ( .IN1(n1734), .IN2(search_data[29]), .S(
        \read_value_mux[30][29] ), .Q(n2646) );
  MUX21X1 U3806 ( .IN1(n1661), .IN2(search_data[0]), .S(
        \read_value_mux[30][0] ), .Q(n2645) );
  MUX21X1 U3807 ( .IN1(n1678), .IN2(search_data[6]), .S(
        \read_value_mux[30][6] ), .Q(n2644) );
  NAND4X0 U3808 ( .IN1(n2647), .IN2(n2646), .IN3(n2645), .IN4(n2644), .QN(
        n2648) );
  NOR4X0 U3809 ( .IN1(n2650), .IN2(n2649), .IN3(n1611), .IN4(n2648), .QN(n2672) );
  MUX21X1 U3810 ( .IN1(n1737), .IN2(search_data[30]), .S(
        \read_value_mux[30][30] ), .Q(n2654) );
  MUX21X1 U3811 ( .IN1(n1694), .IN2(search_data[11]), .S(
        \read_value_mux[30][11] ), .Q(n2653) );
  MUX21X1 U3812 ( .IN1(n1709), .IN2(search_data[17]), .S(
        \read_value_mux[30][17] ), .Q(n2652) );
  MUX21X1 U3813 ( .IN1(n1663), .IN2(search_data[1]), .S(
        \read_value_mux[30][1] ), .Q(n2651) );
  NAND4X0 U3814 ( .IN1(n2654), .IN2(n2653), .IN3(n2652), .IN4(n2651), .QN(
        n2670) );
  MUX21X1 U3815 ( .IN1(n1696), .IN2(search_data[12]), .S(
        \read_value_mux[30][12] ), .Q(n2658) );
  MUX21X1 U3816 ( .IN1(n1672), .IN2(search_data[4]), .S(
        \read_value_mux[30][4] ), .Q(n2657) );
  MUX21X1 U3817 ( .IN1(n1719), .IN2(search_data[21]), .S(
        \read_value_mux[30][21] ), .Q(n2656) );
  MUX21X1 U3818 ( .IN1(n1713), .IN2(search_data[18]), .S(
        \read_value_mux[30][18] ), .Q(n2655) );
  NAND4X0 U3819 ( .IN1(n2658), .IN2(n2657), .IN3(n2656), .IN4(n2655), .QN(
        n2669) );
  MUX21X1 U3820 ( .IN1(n1707), .IN2(search_data[16]), .S(
        \read_value_mux[30][16] ), .Q(n2661) );
  MUX21X1 U3821 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[30][25] ), .Q(n2660) );
  MUX21X1 U3822 ( .IN1(n1731), .IN2(search_data[27]), .S(
        \read_value_mux[30][27] ), .Q(n2659) );
  NAND4X0 U3823 ( .IN1(n2662), .IN2(n2661), .IN3(n2660), .IN4(n2659), .QN(
        n2668) );
  MUX21X1 U3824 ( .IN1(n1692), .IN2(search_data[10]), .S(
        \read_value_mux[30][10] ), .Q(n2666) );
  MUX21X1 U3825 ( .IN1(n1718), .IN2(search_data[20]), .S(
        \read_value_mux[30][20] ), .Q(n2665) );
  MUX21X1 U3826 ( .IN1(n1716), .IN2(search_data[19]), .S(
        \read_value_mux[30][19] ), .Q(n2664) );
  MUX21X1 U3827 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[30][23] ), .Q(n2663) );
  NAND4X0 U3828 ( .IN1(n2666), .IN2(n2665), .IN3(n2664), .IN4(n2663), .QN(
        n2667) );
  NOR4X0 U3829 ( .IN1(n2670), .IN2(n2669), .IN3(n2668), .IN4(n2667), .QN(n2671) );
  NAND4X0 U3830 ( .IN1(n2674), .IN2(n2673), .IN3(n2672), .IN4(n2671), .QN(
        n3076) );
  MUX21X1 U3831 ( .IN1(n1690), .IN2(n1691), .S(\read_value_mux[28][10] ), .Q(
        n2683) );
  MUX21X1 U3832 ( .IN1(search_data[17]), .IN2(n1709), .S(
        \read_value_mux[28][17] ), .Q(n2682) );
  OAI22X1 U3833 ( .IN1(\read_value_mux[28][0] ), .IN2(n1661), .IN3(n1686), 
        .IN4(\read_value_mux[28][8] ), .QN(n2675) );
  AO221X1 U3834 ( .IN1(n1661), .IN2(\read_value_mux[28][0] ), .IN3(n1686), 
        .IN4(\read_value_mux[28][8] ), .IN5(n2675), .Q(n2681) );
  MUX21X1 U3835 ( .IN1(n1719), .IN2(search_data[21]), .S(
        \read_value_mux[28][21] ), .Q(n2679) );
  MUX21X1 U3836 ( .IN1(n1675), .IN2(search_data[5]), .S(
        \read_value_mux[28][5] ), .Q(n2678) );
  MUX21X1 U3837 ( .IN1(n1701), .IN2(search_data[14]), .S(
        \read_value_mux[28][14] ), .Q(n2677) );
  MUX21X1 U3838 ( .IN1(n1728), .IN2(search_data[26]), .S(
        \read_value_mux[28][26] ), .Q(n2676) );
  NAND4X0 U3839 ( .IN1(n2679), .IN2(n2678), .IN3(n2677), .IN4(n2676), .QN(
        n2680) );
  NOR4X0 U3840 ( .IN1(n2683), .IN2(n2682), .IN3(n2681), .IN4(n2680), .QN(n2715) );
  AOI22X1 U3841 ( .IN1(n1683), .IN2(\read_value_mux[28][7] ), .IN3(n1706), 
        .IN4(\read_value_mux[28][15] ), .QN(n2684) );
  OA221X1 U3842 ( .IN1(n1683), .IN2(\read_value_mux[28][7] ), .IN3(n1706), 
        .IN4(\read_value_mux[28][15] ), .IN5(n2684), .Q(n2714) );
  MUX21X1 U3843 ( .IN1(search_data[27]), .IN2(n1730), .S(
        \read_value_mux[28][27] ), .Q(n2691) );
  MUX21X1 U3844 ( .IN1(search_data[25]), .IN2(n1727), .S(
        \read_value_mux[28][25] ), .Q(n2690) );
  MUX21X1 U3845 ( .IN1(n1738), .IN2(search_data[30]), .S(
        \read_value_mux[28][30] ), .Q(n2688) );
  MUX21X1 U3846 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[28][24] ), .Q(n2687) );
  MUX21X1 U3847 ( .IN1(n1734), .IN2(search_data[29]), .S(
        \read_value_mux[28][29] ), .Q(n2686) );
  NAND4X0 U3848 ( .IN1(n2688), .IN2(n2687), .IN3(n2686), .IN4(n2685), .QN(
        n2689) );
  NOR4X0 U3849 ( .IN1(n2691), .IN2(n2690), .IN3(n1611), .IN4(n2689), .QN(n2713) );
  MUX21X1 U3850 ( .IN1(n1672), .IN2(search_data[4]), .S(
        \read_value_mux[28][4] ), .Q(n2695) );
  MUX21X1 U3851 ( .IN1(n1687), .IN2(search_data[9]), .S(
        \read_value_mux[28][9] ), .Q(n2694) );
  MUX21X1 U3852 ( .IN1(n1678), .IN2(search_data[6]), .S(
        \read_value_mux[28][6] ), .Q(n2693) );
  MUX21X1 U3853 ( .IN1(n1696), .IN2(search_data[12]), .S(
        \read_value_mux[28][12] ), .Q(n2692) );
  NAND4X0 U3854 ( .IN1(n2695), .IN2(n2694), .IN3(n2693), .IN4(n2692), .QN(
        n2711) );
  MUX21X1 U3855 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[28][23] ), .Q(n2699) );
  MUX21X1 U3856 ( .IN1(n1663), .IN2(search_data[1]), .S(
        \read_value_mux[28][1] ), .Q(n2698) );
  MUX21X1 U3857 ( .IN1(n1669), .IN2(search_data[3]), .S(
        \read_value_mux[28][3] ), .Q(n2697) );
  MUX21X1 U3858 ( .IN1(n1708), .IN2(search_data[16]), .S(
        \read_value_mux[28][16] ), .Q(n2696) );
  NAND4X0 U3859 ( .IN1(n2699), .IN2(n2698), .IN3(n2697), .IN4(n2696), .QN(
        n2710) );
  MUX21X1 U3860 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[28][28] ), .Q(n2703) );
  MUX21X1 U3861 ( .IN1(n1694), .IN2(search_data[11]), .S(
        \read_value_mux[28][11] ), .Q(n2702) );
  MUX21X1 U3862 ( .IN1(n1722), .IN2(search_data[22]), .S(
        \read_value_mux[28][22] ), .Q(n2701) );
  MUX21X1 U3863 ( .IN1(n1716), .IN2(search_data[19]), .S(
        \read_value_mux[28][19] ), .Q(n2700) );
  NAND4X0 U3864 ( .IN1(n2703), .IN2(n2702), .IN3(n2701), .IN4(n2700), .QN(
        n2709) );
  MUX21X1 U3865 ( .IN1(n1666), .IN2(search_data[2]), .S(
        \read_value_mux[28][2] ), .Q(n2707) );
  MUX21X1 U3866 ( .IN1(n1713), .IN2(search_data[18]), .S(
        \read_value_mux[28][18] ), .Q(n2706) );
  MUX21X1 U3867 ( .IN1(n1741), .IN2(search_data[31]), .S(
        \read_value_mux[28][31] ), .Q(n2705) );
  MUX21X1 U3868 ( .IN1(n1718), .IN2(search_data[20]), .S(
        \read_value_mux[28][20] ), .Q(n2704) );
  NAND4X0 U3869 ( .IN1(n2707), .IN2(n2706), .IN3(n2705), .IN4(n2704), .QN(
        n2708) );
  NOR4X0 U3870 ( .IN1(n2711), .IN2(n2710), .IN3(n2709), .IN4(n2708), .QN(n2712) );
  NAND4X0 U3871 ( .IN1(n2715), .IN2(n2714), .IN3(n2713), .IN4(n2712), .QN(
        n3079) );
  OA221X1 U3872 ( .IN1(n3077), .IN2(n3074), .IN3(n3077), .IN4(n3076), .IN5(
        n3079), .Q(n2755) );
  AOI22X1 U3873 ( .IN1(n1665), .IN2(\read_value_mux[25][1] ), .IN3(n1732), 
        .IN4(\read_value_mux[25][27] ), .QN(n2716) );
  OA221X1 U3874 ( .IN1(n1665), .IN2(\read_value_mux[25][1] ), .IN3(n1732), 
        .IN4(\read_value_mux[25][27] ), .IN5(n2716), .Q(n2721) );
  AOI22X1 U3875 ( .IN1(n1683), .IN2(\read_value_mux[25][7] ), .IN3(n1708), 
        .IN4(\read_value_mux[25][16] ), .QN(n2717) );
  OA221X1 U3876 ( .IN1(n1683), .IN2(\read_value_mux[25][7] ), .IN3(n1708), 
        .IN4(\read_value_mux[25][16] ), .IN5(n2717), .Q(n2720) );
  MUX21X1 U3877 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[25][28] ), .Q(n2719) );
  MUX21X1 U3878 ( .IN1(n1672), .IN2(search_data[4]), .S(
        \read_value_mux[25][4] ), .Q(n2718) );
  NAND4X0 U3879 ( .IN1(n2721), .IN2(n2720), .IN3(n2719), .IN4(n2718), .QN(
        n2754) );
  MUX21X1 U3880 ( .IN1(search_data[20]), .IN2(n1718), .S(
        \read_value_mux[25][20] ), .Q(n2728) );
  MUX21X1 U3881 ( .IN1(search_data[6]), .IN2(n1678), .S(
        \read_value_mux[25][6] ), .Q(n2727) );
  MUX21X1 U3882 ( .IN1(n1719), .IN2(search_data[21]), .S(
        \read_value_mux[25][21] ), .Q(n2725) );
  MUX21X1 U3883 ( .IN1(n1684), .IN2(search_data[8]), .S(
        \read_value_mux[25][8] ), .Q(n2724) );
  MUX21X1 U3884 ( .IN1(n1709), .IN2(search_data[17]), .S(
        \read_value_mux[25][17] ), .Q(n2723) );
  MUX21X1 U3885 ( .IN1(n1666), .IN2(search_data[2]), .S(
        \read_value_mux[25][2] ), .Q(n2722) );
  NAND4X0 U3886 ( .IN1(n2725), .IN2(n2724), .IN3(n2723), .IN4(n2722), .QN(
        n2726) );
  NOR4X0 U3887 ( .IN1(n2728), .IN2(n2727), .IN3(n1611), .IN4(n2726), .QN(n2752) );
  MUX21X1 U3888 ( .IN1(n1713), .IN2(search_data[18]), .S(
        \read_value_mux[25][18] ), .Q(n2732) );
  MUX21X1 U3889 ( .IN1(n1705), .IN2(n1704), .S(\read_value_mux[25][15] ), .Q(
        n2731) );
  MUX21X1 U3890 ( .IN1(n1693), .IN2(search_data[11]), .S(
        \read_value_mux[25][11] ), .Q(n2730) );
  MUX21X1 U3891 ( .IN1(n1687), .IN2(search_data[9]), .S(
        \read_value_mux[25][9] ), .Q(n2729) );
  NAND4X0 U3892 ( .IN1(n2732), .IN2(n2731), .IN3(n2730), .IN4(n2729), .QN(
        n2748) );
  MUX21X1 U3893 ( .IN1(n1722), .IN2(search_data[22]), .S(
        \read_value_mux[25][22] ), .Q(n2736) );
  MUX21X1 U3894 ( .IN1(n1698), .IN2(search_data[13]), .S(
        \read_value_mux[25][13] ), .Q(n2735) );
  MUX21X1 U3895 ( .IN1(n1737), .IN2(search_data[30]), .S(
        \read_value_mux[25][30] ), .Q(n2733) );
  NAND4X0 U3896 ( .IN1(n2736), .IN2(n2735), .IN3(n2734), .IN4(n2733), .QN(
        n2747) );
  MUX21X1 U3897 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[25][23] ), .Q(n2740) );
  MUX21X1 U3898 ( .IN1(n1740), .IN2(search_data[31]), .S(
        \read_value_mux[25][31] ), .Q(n2739) );
  MUX21X1 U3899 ( .IN1(n1697), .IN2(search_data[12]), .S(
        \read_value_mux[25][12] ), .Q(n2738) );
  MUX21X1 U3900 ( .IN1(n1701), .IN2(search_data[14]), .S(
        \read_value_mux[25][14] ), .Q(n2737) );
  NAND4X0 U3901 ( .IN1(n2740), .IN2(n2739), .IN3(n2738), .IN4(n2737), .QN(
        n2746) );
  MUX21X1 U3902 ( .IN1(n1717), .IN2(search_data[19]), .S(
        \read_value_mux[25][19] ), .Q(n2744) );
  MUX21X1 U3903 ( .IN1(n1669), .IN2(search_data[3]), .S(
        \read_value_mux[25][3] ), .Q(n2742) );
  MUX21X1 U3904 ( .IN1(n1734), .IN2(search_data[29]), .S(
        \read_value_mux[25][29] ), .Q(n2741) );
  NAND4X0 U3905 ( .IN1(n2744), .IN2(n2743), .IN3(n2742), .IN4(n2741), .QN(
        n2745) );
  NOR4X0 U3906 ( .IN1(n2748), .IN2(n2747), .IN3(n2746), .IN4(n2745), .QN(n2751) );
  MUX21X1 U3907 ( .IN1(n1675), .IN2(search_data[5]), .S(
        \read_value_mux[25][5] ), .Q(n2750) );
  MUX21X1 U3908 ( .IN1(n1661), .IN2(search_data[0]), .S(
        \read_value_mux[25][0] ), .Q(n2749) );
  NAND4X0 U3909 ( .IN1(n2752), .IN2(n2751), .IN3(n2750), .IN4(n2749), .QN(
        n2753) );
  AO221X1 U3910 ( .IN1(n3071), .IN2(n3072), .IN3(n3071), .IN4(n2755), .IN5(
        n3080), .Q(n2797) );
  MUX21X1 U3911 ( .IN1(search_data[1]), .IN2(n1663), .S(
        \read_value_mux[22][1] ), .Q(n2764) );
  MUX21X1 U3912 ( .IN1(search_data[3]), .IN2(n1669), .S(
        \read_value_mux[22][3] ), .Q(n2763) );
  OAI22X1 U3913 ( .IN1(n1661), .IN2(\read_value_mux[22][0] ), .IN3(n1674), 
        .IN4(\read_value_mux[22][4] ), .QN(n2756) );
  AO221X1 U3914 ( .IN1(n1661), .IN2(\read_value_mux[22][0] ), .IN3(
        \read_value_mux[22][4] ), .IN4(n1674), .IN5(n2756), .Q(n2762) );
  MUX21X1 U3915 ( .IN1(n1728), .IN2(search_data[26]), .S(
        \read_value_mux[22][26] ), .Q(n2760) );
  MUX21X1 U3916 ( .IN1(n1698), .IN2(search_data[13]), .S(
        \read_value_mux[22][13] ), .Q(n2759) );
  MUX21X1 U3917 ( .IN1(n1693), .IN2(search_data[11]), .S(
        \read_value_mux[22][11] ), .Q(n2758) );
  MUX21X1 U3918 ( .IN1(n1740), .IN2(search_data[31]), .S(
        \read_value_mux[22][31] ), .Q(n2757) );
  NAND4X0 U3919 ( .IN1(n2760), .IN2(n2759), .IN3(n2758), .IN4(n2757), .QN(
        n2761) );
  NOR4X0 U3920 ( .IN1(n2764), .IN2(n2763), .IN3(n2762), .IN4(n2761), .QN(n2796) );
  AOI22X1 U3921 ( .IN1(n1691), .IN2(\read_value_mux[22][10] ), .IN3(n1732), 
        .IN4(\read_value_mux[22][27] ), .QN(n2765) );
  OA221X1 U3922 ( .IN1(n1691), .IN2(\read_value_mux[22][10] ), .IN3(n1732), 
        .IN4(\read_value_mux[22][27] ), .IN5(n2765), .Q(n2795) );
  MUX21X1 U3923 ( .IN1(search_data[19]), .IN2(n1717), .S(
        \read_value_mux[22][19] ), .Q(n2772) );
  MUX21X1 U3924 ( .IN1(search_data[20]), .IN2(n1718), .S(
        \read_value_mux[22][20] ), .Q(n2771) );
  MUX21X1 U3925 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[22][28] ), .Q(n2769) );
  MUX21X1 U3926 ( .IN1(n1701), .IN2(search_data[14]), .S(
        \read_value_mux[22][14] ), .Q(n2768) );
  MUX21X1 U3927 ( .IN1(n1684), .IN2(search_data[8]), .S(
        \read_value_mux[22][8] ), .Q(n2767) );
  MUX21X1 U3928 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[22][25] ), .Q(n2766) );
  NAND4X0 U3929 ( .IN1(n2769), .IN2(n2768), .IN3(n2767), .IN4(n2766), .QN(
        n2770) );
  NOR4X0 U3930 ( .IN1(n2772), .IN2(n2771), .IN3(n1611), .IN4(n2770), .QN(n2794) );
  MUX21X1 U3931 ( .IN1(n1666), .IN2(search_data[2]), .S(
        \read_value_mux[22][2] ), .Q(n2776) );
  MUX21X1 U3932 ( .IN1(n1697), .IN2(search_data[12]), .S(
        \read_value_mux[22][12] ), .Q(n2775) );
  MUX21X1 U3933 ( .IN1(n1722), .IN2(search_data[22]), .S(
        \read_value_mux[22][22] ), .Q(n2774) );
  MUX21X1 U3934 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[22][23] ), .Q(n2773) );
  NAND4X0 U3935 ( .IN1(n2776), .IN2(n2775), .IN3(n2774), .IN4(n2773), .QN(
        n2792) );
  MUX21X1 U3936 ( .IN1(n1705), .IN2(n1704), .S(\read_value_mux[22][15] ), .Q(
        n2780) );
  MUX21X1 U3937 ( .IN1(n1707), .IN2(search_data[16]), .S(
        \read_value_mux[22][16] ), .Q(n2779) );
  MUX21X1 U3938 ( .IN1(n1675), .IN2(search_data[5]), .S(
        \read_value_mux[22][5] ), .Q(n2778) );
  MUX21X1 U3939 ( .IN1(n1737), .IN2(search_data[30]), .S(
        \read_value_mux[22][30] ), .Q(n2777) );
  NAND4X0 U3940 ( .IN1(n2780), .IN2(n2779), .IN3(n2778), .IN4(n2777), .QN(
        n2791) );
  MUX21X1 U3941 ( .IN1(n1709), .IN2(search_data[17]), .S(
        \read_value_mux[22][17] ), .Q(n2784) );
  MUX21X1 U3942 ( .IN1(n1720), .IN2(search_data[21]), .S(
        \read_value_mux[22][21] ), .Q(n2783) );
  MUX21X1 U3943 ( .IN1(n1678), .IN2(search_data[6]), .S(
        \read_value_mux[22][6] ), .Q(n2782) );
  MUX21X1 U3944 ( .IN1(n1681), .IN2(search_data[7]), .S(
        \read_value_mux[22][7] ), .Q(n2781) );
  NAND4X0 U3945 ( .IN1(n2784), .IN2(n2783), .IN3(n2782), .IN4(n2781), .QN(
        n2790) );
  MUX21X1 U3946 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[22][24] ), .Q(n2788) );
  MUX21X1 U3947 ( .IN1(n1734), .IN2(search_data[29]), .S(
        \read_value_mux[22][29] ), .Q(n2787) );
  MUX21X1 U3948 ( .IN1(n1714), .IN2(search_data[18]), .S(
        \read_value_mux[22][18] ), .Q(n2786) );
  MUX21X1 U3949 ( .IN1(n1687), .IN2(search_data[9]), .S(
        \read_value_mux[22][9] ), .Q(n2785) );
  NAND4X0 U3950 ( .IN1(n2788), .IN2(n2787), .IN3(n2786), .IN4(n2785), .QN(
        n2789) );
  NOR4X0 U3951 ( .IN1(n2792), .IN2(n2791), .IN3(n2790), .IN4(n2789), .QN(n2793) );
  NAND4X0 U3952 ( .IN1(n2796), .IN2(n2795), .IN3(n2794), .IN4(n2793), .QN(
        n3070) );
  OA221X1 U3953 ( .IN1(n3068), .IN2(n3111), .IN3(n3068), .IN4(n2797), .IN5(
        n3070), .Q(n2839) );
  MUX21X1 U3954 ( .IN1(search_data[27]), .IN2(n1730), .S(
        \read_value_mux[19][27] ), .Q(n2838) );
  MUX21X1 U3955 ( .IN1(search_data[30]), .IN2(n1737), .S(
        \read_value_mux[19][30] ), .Q(n2837) );
  AOI22X1 U3956 ( .IN1(n1697), .IN2(\read_value_mux[19][12] ), .IN3(n1703), 
        .IN4(\read_value_mux[19][14] ), .QN(n2798) );
  OA221X1 U3957 ( .IN1(n1697), .IN2(\read_value_mux[19][12] ), .IN3(n1703), 
        .IN4(\read_value_mux[19][14] ), .IN5(n2798), .Q(n2803) );
  AOI22X1 U3958 ( .IN1(n1668), .IN2(\read_value_mux[19][2] ), .IN3(n1718), 
        .IN4(\read_value_mux[19][20] ), .QN(n2799) );
  OA221X1 U3959 ( .IN1(n1668), .IN2(\read_value_mux[19][2] ), .IN3(n1718), 
        .IN4(\read_value_mux[19][20] ), .IN5(n2799), .Q(n2802) );
  MUX21X1 U3960 ( .IN1(n1693), .IN2(search_data[11]), .S(
        \read_value_mux[19][11] ), .Q(n2801) );
  MUX21X1 U3961 ( .IN1(n1698), .IN2(search_data[13]), .S(
        \read_value_mux[19][13] ), .Q(n2800) );
  NAND4X0 U3962 ( .IN1(n2803), .IN2(n2802), .IN3(n2801), .IN4(n2800), .QN(
        n2836) );
  MUX21X1 U3963 ( .IN1(search_data[24]), .IN2(n1726), .S(
        \read_value_mux[19][24] ), .Q(n2810) );
  MUX21X1 U3964 ( .IN1(search_data[31]), .IN2(n1740), .S(
        \read_value_mux[19][31] ), .Q(n2809) );
  MUX21X1 U3965 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[19][23] ), .Q(n2807) );
  MUX21X1 U3966 ( .IN1(n1713), .IN2(search_data[18]), .S(
        \read_value_mux[19][18] ), .Q(n2806) );
  MUX21X1 U3967 ( .IN1(n1681), .IN2(search_data[7]), .S(
        \read_value_mux[19][7] ), .Q(n2805) );
  MUX21X1 U3968 ( .IN1(n1663), .IN2(search_data[1]), .S(
        \read_value_mux[19][1] ), .Q(n2804) );
  NAND4X0 U3969 ( .IN1(n2807), .IN2(n2806), .IN3(n2805), .IN4(n2804), .QN(
        n2808) );
  NOR4X0 U3970 ( .IN1(n2810), .IN2(n2809), .IN3(n1611), .IN4(n2808), .QN(n2834) );
  MUX21X1 U3971 ( .IN1(n1728), .IN2(search_data[26]), .S(
        \read_value_mux[19][26] ), .Q(n2814) );
  MUX21X1 U3972 ( .IN1(n1691), .IN2(search_data[10]), .S(
        \read_value_mux[19][10] ), .Q(n2813) );
  MUX21X1 U3973 ( .IN1(n1709), .IN2(search_data[17]), .S(
        \read_value_mux[19][17] ), .Q(n2812) );
  MUX21X1 U3974 ( .IN1(n1660), .IN2(search_data[0]), .S(
        \read_value_mux[19][0] ), .Q(n2811) );
  NAND4X0 U3975 ( .IN1(n2814), .IN2(n2813), .IN3(n2812), .IN4(n2811), .QN(
        n2830) );
  MUX21X1 U3976 ( .IN1(n1672), .IN2(search_data[4]), .S(
        \read_value_mux[19][4] ), .Q(n2818) );
  MUX21X1 U3977 ( .IN1(n1687), .IN2(search_data[9]), .S(
        \read_value_mux[19][9] ), .Q(n2817) );
  MUX21X1 U3978 ( .IN1(n1719), .IN2(search_data[21]), .S(
        \read_value_mux[19][21] ), .Q(n2816) );
  MUX21X1 U3979 ( .IN1(n1678), .IN2(search_data[6]), .S(
        \read_value_mux[19][6] ), .Q(n2815) );
  NAND4X0 U3980 ( .IN1(n2818), .IN2(n2817), .IN3(n2816), .IN4(n2815), .QN(
        n2829) );
  MUX21X1 U3981 ( .IN1(n1716), .IN2(search_data[19]), .S(
        \read_value_mux[19][19] ), .Q(n2822) );
  MUX21X1 U3982 ( .IN1(n1669), .IN2(search_data[3]), .S(
        \read_value_mux[19][3] ), .Q(n2821) );
  MUX21X1 U3983 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[19][28] ), .Q(n2820) );
  MUX21X1 U3984 ( .IN1(n1675), .IN2(search_data[5]), .S(
        \read_value_mux[19][5] ), .Q(n2819) );
  NAND4X0 U3985 ( .IN1(n2822), .IN2(n2821), .IN3(n2820), .IN4(n2819), .QN(
        n2828) );
  MUX21X1 U3986 ( .IN1(n1734), .IN2(search_data[29]), .S(
        \read_value_mux[19][29] ), .Q(n2826) );
  MUX21X1 U3987 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[19][25] ), .Q(n2825) );
  MUX21X1 U3988 ( .IN1(n1708), .IN2(search_data[16]), .S(
        \read_value_mux[19][16] ), .Q(n2824) );
  MUX21X1 U3989 ( .IN1(n1684), .IN2(search_data[8]), .S(
        \read_value_mux[19][8] ), .Q(n2823) );
  NAND4X0 U3990 ( .IN1(n2826), .IN2(n2825), .IN3(n2824), .IN4(n2823), .QN(
        n2827) );
  NOR4X0 U3991 ( .IN1(n2830), .IN2(n2829), .IN3(n2828), .IN4(n2827), .QN(n2833) );
  MUX21X1 U3992 ( .IN1(n1722), .IN2(search_data[22]), .S(
        \read_value_mux[19][22] ), .Q(n2832) );
  MUX21X1 U3993 ( .IN1(n1705), .IN2(n1704), .S(\read_value_mux[19][15] ), .Q(
        n2831) );
  NAND4X0 U3994 ( .IN1(n2834), .IN2(n2833), .IN3(n2832), .IN4(n2831), .QN(
        n2835) );
  NOR4X0 U3995 ( .IN1(n2838), .IN2(n2837), .IN3(n2836), .IN4(n2835), .QN(n3083) );
  AO221X1 U3996 ( .IN1(n3067), .IN2(n3065), .IN3(n3067), .IN4(n2839), .IN5(
        n3083), .Q(n2840) );
  MUX21X1 U3997 ( .IN1(search_data[18]), .IN2(n1712), .S(
        \read_value_mux[11][18] ), .Q(n2881) );
  MUX21X1 U3998 ( .IN1(search_data[2]), .IN2(n1666), .S(
        \read_value_mux[11][2] ), .Q(n2880) );
  AOI22X1 U3999 ( .IN1(n1686), .IN2(\read_value_mux[11][8] ), .IN3(n1703), 
        .IN4(\read_value_mux[11][14] ), .QN(n2841) );
  OA221X1 U4000 ( .IN1(n1686), .IN2(\read_value_mux[11][8] ), .IN3(n1703), 
        .IN4(\read_value_mux[11][14] ), .IN5(n2841), .Q(n2846) );
  AOI22X1 U4001 ( .IN1(n1727), .IN2(\read_value_mux[11][25] ), .IN3(n1677), 
        .IN4(\read_value_mux[11][5] ), .QN(n2842) );
  OA221X1 U4002 ( .IN1(n1727), .IN2(\read_value_mux[11][25] ), .IN3(n1677), 
        .IN4(\read_value_mux[11][5] ), .IN5(n2842), .Q(n2845) );
  MUX21X1 U4003 ( .IN1(n1722), .IN2(search_data[22]), .S(
        \read_value_mux[11][22] ), .Q(n2844) );
  MUX21X1 U4004 ( .IN1(n1687), .IN2(search_data[9]), .S(
        \read_value_mux[11][9] ), .Q(n2843) );
  NAND4X0 U4005 ( .IN1(n2846), .IN2(n2845), .IN3(n2844), .IN4(n2843), .QN(
        n2879) );
  MUX21X1 U4006 ( .IN1(search_data[19]), .IN2(n1717), .S(
        \read_value_mux[11][19] ), .Q(n2853) );
  MUX21X1 U4007 ( .IN1(search_data[21]), .IN2(n1719), .S(
        \read_value_mux[11][21] ), .Q(n2852) );
  MUX21X1 U4008 ( .IN1(n1696), .IN2(search_data[12]), .S(
        \read_value_mux[11][12] ), .Q(n2850) );
  MUX21X1 U4009 ( .IN1(n1707), .IN2(search_data[16]), .S(
        \read_value_mux[11][16] ), .Q(n2849) );
  MUX21X1 U4010 ( .IN1(n1705), .IN2(n1704), .S(\read_value_mux[11][15] ), .Q(
        n2848) );
  MUX21X1 U4011 ( .IN1(n1698), .IN2(search_data[13]), .S(
        \read_value_mux[11][13] ), .Q(n2847) );
  NAND4X0 U4012 ( .IN1(n2850), .IN2(n2849), .IN3(n2848), .IN4(n2847), .QN(
        n2851) );
  NOR4X0 U4013 ( .IN1(n2853), .IN2(n2852), .IN3(n1611), .IN4(n2851), .QN(n2877) );
  MUX21X1 U4014 ( .IN1(n1681), .IN2(search_data[7]), .S(
        \read_value_mux[11][7] ), .Q(n2857) );
  MUX21X1 U4015 ( .IN1(n1734), .IN2(search_data[29]), .S(
        \read_value_mux[11][29] ), .Q(n2856) );
  MUX21X1 U4016 ( .IN1(n1740), .IN2(search_data[31]), .S(
        \read_value_mux[11][31] ), .Q(n2855) );
  MUX21X1 U4017 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[11][24] ), .Q(n2854) );
  NAND4X0 U4018 ( .IN1(n2857), .IN2(n2856), .IN3(n2855), .IN4(n2854), .QN(
        n2873) );
  MUX21X1 U4019 ( .IN1(n1709), .IN2(search_data[17]), .S(
        \read_value_mux[11][17] ), .Q(n2861) );
  MUX21X1 U4020 ( .IN1(n1693), .IN2(search_data[11]), .S(
        \read_value_mux[11][11] ), .Q(n2860) );
  MUX21X1 U4021 ( .IN1(n1691), .IN2(search_data[10]), .S(
        \read_value_mux[11][10] ), .Q(n2859) );
  MUX21X1 U4022 ( .IN1(n1728), .IN2(search_data[26]), .S(
        \read_value_mux[11][26] ), .Q(n2858) );
  NAND4X0 U4023 ( .IN1(n2861), .IN2(n2860), .IN3(n2859), .IN4(n2858), .QN(
        n2872) );
  MUX21X1 U4024 ( .IN1(n1664), .IN2(search_data[1]), .S(
        \read_value_mux[11][1] ), .Q(n2865) );
  MUX21X1 U4025 ( .IN1(n1678), .IN2(search_data[6]), .S(
        \read_value_mux[11][6] ), .Q(n2864) );
  MUX21X1 U4026 ( .IN1(n1660), .IN2(search_data[0]), .S(
        \read_value_mux[11][0] ), .Q(n2863) );
  MUX21X1 U4027 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[11][28] ), .Q(n2862) );
  NAND4X0 U4028 ( .IN1(n2865), .IN2(n2864), .IN3(n2863), .IN4(n2862), .QN(
        n2871) );
  MUX21X1 U4029 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[11][23] ), .Q(n2869) );
  MUX21X1 U4030 ( .IN1(n1669), .IN2(search_data[3]), .S(
        \read_value_mux[11][3] ), .Q(n2868) );
  MUX21X1 U4031 ( .IN1(n1718), .IN2(search_data[20]), .S(
        \read_value_mux[11][20] ), .Q(n2867) );
  MUX21X1 U4032 ( .IN1(n1731), .IN2(search_data[27]), .S(
        \read_value_mux[11][27] ), .Q(n2866) );
  NAND4X0 U4033 ( .IN1(n2869), .IN2(n2868), .IN3(n2867), .IN4(n2866), .QN(
        n2870) );
  NOR4X0 U4034 ( .IN1(n2873), .IN2(n2872), .IN3(n2871), .IN4(n2870), .QN(n2876) );
  MUX21X1 U4035 ( .IN1(n1672), .IN2(search_data[4]), .S(
        \read_value_mux[11][4] ), .Q(n2875) );
  MUX21X1 U4036 ( .IN1(n1737), .IN2(search_data[30]), .S(
        \read_value_mux[11][30] ), .Q(n2874) );
  NAND4X0 U4037 ( .IN1(n2877), .IN2(n2876), .IN3(n2875), .IN4(n2874), .QN(
        n2878) );
  NOR4X0 U4038 ( .IN1(n2881), .IN2(n2880), .IN3(n2879), .IN4(n2878), .QN(n3063) );
  MUX21X1 U4039 ( .IN1(search_data[28]), .IN2(n1733), .S(
        \read_value_mux[15][28] ), .Q(n2922) );
  MUX21X1 U4040 ( .IN1(search_data[6]), .IN2(n1678), .S(
        \read_value_mux[15][6] ), .Q(n2921) );
  AOI22X1 U4041 ( .IN1(n1726), .IN2(\read_value_mux[15][24] ), .IN3(n1697), 
        .IN4(\read_value_mux[15][12] ), .QN(n2882) );
  OA221X1 U4042 ( .IN1(n1726), .IN2(\read_value_mux[15][24] ), .IN3(n1697), 
        .IN4(\read_value_mux[15][12] ), .IN5(n2882), .Q(n2887) );
  AOI22X1 U4043 ( .IN1(n1661), .IN2(\read_value_mux[15][0] ), .IN3(n1732), 
        .IN4(\read_value_mux[15][27] ), .QN(n2883) );
  OA221X1 U4044 ( .IN1(n1661), .IN2(\read_value_mux[15][0] ), .IN3(n1732), 
        .IN4(\read_value_mux[15][27] ), .IN5(n2883), .Q(n2886) );
  MUX21X1 U4045 ( .IN1(n1740), .IN2(search_data[31]), .S(
        \read_value_mux[15][31] ), .Q(n2885) );
  MUX21X1 U4046 ( .IN1(n1715), .IN2(search_data[19]), .S(
        \read_value_mux[15][19] ), .Q(n2884) );
  NAND4X0 U4047 ( .IN1(n2887), .IN2(n2886), .IN3(n2885), .IN4(n2884), .QN(
        n2920) );
  MUX21X1 U4048 ( .IN1(search_data[7]), .IN2(n1681), .S(
        \read_value_mux[15][7] ), .Q(n2894) );
  MUX21X1 U4049 ( .IN1(search_data[25]), .IN2(n1727), .S(
        \read_value_mux[15][25] ), .Q(n2893) );
  MUX21X1 U4050 ( .IN1(n1663), .IN2(search_data[1]), .S(
        \read_value_mux[15][1] ), .Q(n2891) );
  MUX21X1 U4051 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[15][23] ), .Q(n2890) );
  MUX21X1 U4052 ( .IN1(n1705), .IN2(n1704), .S(\read_value_mux[15][15] ), .Q(
        n2889) );
  MUX21X1 U4053 ( .IN1(n1687), .IN2(search_data[9]), .S(
        \read_value_mux[15][9] ), .Q(n2888) );
  NAND4X0 U4054 ( .IN1(n2891), .IN2(n2890), .IN3(n2889), .IN4(n2888), .QN(
        n2892) );
  NOR4X0 U4055 ( .IN1(n2894), .IN2(n2893), .IN3(n1611), .IN4(n2892), .QN(n2918) );
  MUX21X1 U4056 ( .IN1(n1693), .IN2(search_data[11]), .S(
        \read_value_mux[15][11] ), .Q(n2898) );
  MUX21X1 U4057 ( .IN1(n1698), .IN2(search_data[13]), .S(
        \read_value_mux[15][13] ), .Q(n2897) );
  MUX21X1 U4058 ( .IN1(n1666), .IN2(search_data[2]), .S(
        \read_value_mux[15][2] ), .Q(n2896) );
  MUX21X1 U4059 ( .IN1(n1701), .IN2(search_data[14]), .S(
        \read_value_mux[15][14] ), .Q(n2895) );
  NAND4X0 U4060 ( .IN1(n2898), .IN2(n2897), .IN3(n2896), .IN4(n2895), .QN(
        n2914) );
  MUX21X1 U4061 ( .IN1(n1691), .IN2(search_data[10]), .S(
        \read_value_mux[15][10] ), .Q(n2902) );
  MUX21X1 U4062 ( .IN1(n1719), .IN2(search_data[21]), .S(
        \read_value_mux[15][21] ), .Q(n2901) );
  MUX21X1 U4063 ( .IN1(n1729), .IN2(search_data[26]), .S(
        \read_value_mux[15][26] ), .Q(n2900) );
  MUX21X1 U4064 ( .IN1(n1718), .IN2(search_data[20]), .S(
        \read_value_mux[15][20] ), .Q(n2899) );
  NAND4X0 U4065 ( .IN1(n2902), .IN2(n2901), .IN3(n2900), .IN4(n2899), .QN(
        n2913) );
  MUX21X1 U4066 ( .IN1(n1709), .IN2(search_data[17]), .S(
        \read_value_mux[15][17] ), .Q(n2906) );
  MUX21X1 U4067 ( .IN1(n1684), .IN2(search_data[8]), .S(
        \read_value_mux[15][8] ), .Q(n2905) );
  MUX21X1 U4068 ( .IN1(n1722), .IN2(search_data[22]), .S(
        \read_value_mux[15][22] ), .Q(n2904) );
  MUX21X1 U4069 ( .IN1(n1734), .IN2(search_data[29]), .S(
        \read_value_mux[15][29] ), .Q(n2903) );
  NAND4X0 U4070 ( .IN1(n2906), .IN2(n2905), .IN3(n2904), .IN4(n2903), .QN(
        n2912) );
  MUX21X1 U4071 ( .IN1(n1708), .IN2(search_data[16]), .S(
        \read_value_mux[15][16] ), .Q(n2910) );
  MUX21X1 U4072 ( .IN1(n1712), .IN2(search_data[18]), .S(
        \read_value_mux[15][18] ), .Q(n2909) );
  MUX21X1 U4073 ( .IN1(n1672), .IN2(search_data[4]), .S(
        \read_value_mux[15][4] ), .Q(n2908) );
  MUX21X1 U4074 ( .IN1(n1737), .IN2(search_data[30]), .S(
        \read_value_mux[15][30] ), .Q(n2907) );
  NAND4X0 U4075 ( .IN1(n2910), .IN2(n2909), .IN3(n2908), .IN4(n2907), .QN(
        n2911) );
  NOR4X0 U4076 ( .IN1(n2914), .IN2(n2913), .IN3(n2912), .IN4(n2911), .QN(n2917) );
  MUX21X1 U4077 ( .IN1(n1675), .IN2(search_data[5]), .S(
        \read_value_mux[15][5] ), .Q(n2916) );
  MUX21X1 U4078 ( .IN1(n1669), .IN2(search_data[3]), .S(
        \read_value_mux[15][3] ), .Q(n2915) );
  NAND4X0 U4079 ( .IN1(n2918), .IN2(n2917), .IN3(n2916), .IN4(n2915), .QN(
        n2919) );
  NOR4X0 U4080 ( .IN1(n2922), .IN2(n2921), .IN3(n2920), .IN4(n2919), .QN(n3089) );
  INVX0 U4081 ( .INP(n2923), .ZN(n2965) );
  MUX21X1 U4082 ( .IN1(search_data[24]), .IN2(n1726), .S(
        \read_value_mux[13][24] ), .Q(n2964) );
  MUX21X1 U4083 ( .IN1(search_data[30]), .IN2(n1737), .S(
        \read_value_mux[13][30] ), .Q(n2963) );
  AOI22X1 U4084 ( .IN1(n1683), .IN2(\read_value_mux[13][7] ), .IN3(n1718), 
        .IN4(\read_value_mux[13][20] ), .QN(n2924) );
  OA221X1 U4085 ( .IN1(n1683), .IN2(\read_value_mux[13][7] ), .IN3(n1718), 
        .IN4(\read_value_mux[13][20] ), .IN5(n2924), .Q(n2929) );
  AOI22X1 U4086 ( .IN1(n1686), .IN2(\read_value_mux[13][8] ), .IN3(n1721), 
        .IN4(\read_value_mux[13][21] ), .QN(n2925) );
  OA221X1 U4087 ( .IN1(n1686), .IN2(\read_value_mux[13][8] ), .IN3(n1721), 
        .IN4(\read_value_mux[13][21] ), .IN5(n2925), .Q(n2928) );
  MUX21X1 U4088 ( .IN1(n1730), .IN2(search_data[27]), .S(
        \read_value_mux[13][27] ), .Q(n2927) );
  MUX21X1 U4089 ( .IN1(n1740), .IN2(search_data[31]), .S(
        \read_value_mux[13][31] ), .Q(n2926) );
  NAND4X0 U4090 ( .IN1(n2929), .IN2(n2928), .IN3(n2927), .IN4(n2926), .QN(
        n2962) );
  MUX21X1 U4091 ( .IN1(search_data[1]), .IN2(n1663), .S(
        \read_value_mux[13][1] ), .Q(n2936) );
  MUX21X1 U4092 ( .IN1(search_data[2]), .IN2(n1666), .S(
        \read_value_mux[13][2] ), .Q(n2935) );
  MUX21X1 U4093 ( .IN1(n1693), .IN2(search_data[11]), .S(
        \read_value_mux[13][11] ), .Q(n2933) );
  MUX21X1 U4094 ( .IN1(n1716), .IN2(search_data[19]), .S(
        \read_value_mux[13][19] ), .Q(n2932) );
  MUX21X1 U4095 ( .IN1(n1698), .IN2(search_data[13]), .S(
        \read_value_mux[13][13] ), .Q(n2931) );
  MUX21X1 U4096 ( .IN1(n1691), .IN2(search_data[10]), .S(
        \read_value_mux[13][10] ), .Q(n2930) );
  NAND4X0 U4097 ( .IN1(n2933), .IN2(n2932), .IN3(n2931), .IN4(n2930), .QN(
        n2934) );
  NOR4X0 U4098 ( .IN1(n2936), .IN2(n2935), .IN3(n1611), .IN4(n2934), .QN(n2960) );
  MUX21X1 U4099 ( .IN1(n1696), .IN2(search_data[12]), .S(
        \read_value_mux[13][12] ), .Q(n2940) );
  MUX21X1 U4100 ( .IN1(n1672), .IN2(search_data[4]), .S(
        \read_value_mux[13][4] ), .Q(n2939) );
  MUX21X1 U4101 ( .IN1(n1669), .IN2(search_data[3]), .S(
        \read_value_mux[13][3] ), .Q(n2938) );
  MUX21X1 U4102 ( .IN1(n1660), .IN2(search_data[0]), .S(
        \read_value_mux[13][0] ), .Q(n2937) );
  NAND4X0 U4103 ( .IN1(n2940), .IN2(n2939), .IN3(n2938), .IN4(n2937), .QN(
        n2956) );
  MUX21X1 U4104 ( .IN1(n1722), .IN2(search_data[22]), .S(
        \read_value_mux[13][22] ), .Q(n2944) );
  MUX21X1 U4105 ( .IN1(n1675), .IN2(search_data[5]), .S(
        \read_value_mux[13][5] ), .Q(n2943) );
  MUX21X1 U4106 ( .IN1(n1705), .IN2(n1704), .S(\read_value_mux[13][15] ), .Q(
        n2942) );
  MUX21X1 U4107 ( .IN1(n1728), .IN2(search_data[26]), .S(
        \read_value_mux[13][26] ), .Q(n2941) );
  NAND4X0 U4108 ( .IN1(n2944), .IN2(n2943), .IN3(n2942), .IN4(n2941), .QN(
        n2955) );
  MUX21X1 U4109 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[13][28] ), .Q(n2948) );
  MUX21X1 U4110 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[13][25] ), .Q(n2947) );
  MUX21X1 U4111 ( .IN1(n1687), .IN2(search_data[9]), .S(
        \read_value_mux[13][9] ), .Q(n2946) );
  MUX21X1 U4112 ( .IN1(n1713), .IN2(search_data[18]), .S(
        \read_value_mux[13][18] ), .Q(n2945) );
  NAND4X0 U4113 ( .IN1(n2948), .IN2(n2947), .IN3(n2946), .IN4(n2945), .QN(
        n2954) );
  MUX21X1 U4114 ( .IN1(n1708), .IN2(search_data[16]), .S(
        \read_value_mux[13][16] ), .Q(n2952) );
  MUX21X1 U4115 ( .IN1(n1701), .IN2(search_data[14]), .S(
        \read_value_mux[13][14] ), .Q(n2951) );
  MUX21X1 U4116 ( .IN1(n1678), .IN2(search_data[6]), .S(
        \read_value_mux[13][6] ), .Q(n2950) );
  MUX21X1 U4117 ( .IN1(n1734), .IN2(search_data[29]), .S(
        \read_value_mux[13][29] ), .Q(n2949) );
  NAND4X0 U4118 ( .IN1(n2952), .IN2(n2951), .IN3(n2950), .IN4(n2949), .QN(
        n2953) );
  NOR4X0 U4119 ( .IN1(n2956), .IN2(n2955), .IN3(n2954), .IN4(n2953), .QN(n2959) );
  MUX21X1 U4120 ( .IN1(n1710), .IN2(search_data[17]), .S(
        \read_value_mux[13][17] ), .Q(n2958) );
  MUX21X1 U4121 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[13][23] ), .Q(n2957) );
  NAND4X0 U4122 ( .IN1(n2960), .IN2(n2959), .IN3(n2958), .IN4(n2957), .QN(
        n2961) );
  NOR4X0 U4123 ( .IN1(n2964), .IN2(n2963), .IN3(n2962), .IN4(n2961), .QN(n3093) );
  AO22X1 U4124 ( .IN1(n3089), .IN2(n2965), .IN3(n3093), .IN4(n3123), .Q(n2966)
         );
  NOR2X0 U4125 ( .IN1(n3063), .IN2(n2966), .QN(n3010) );
  MUX21X1 U4126 ( .IN1(search_data[3]), .IN2(n1669), .S(
        \read_value_mux[17][3] ), .Q(n2975) );
  MUX21X1 U4127 ( .IN1(search_data[17]), .IN2(n1709), .S(
        \read_value_mux[17][17] ), .Q(n2974) );
  OAI22X1 U4128 ( .IN1(n1697), .IN2(\read_value_mux[17][12] ), .IN3(n1721), 
        .IN4(\read_value_mux[17][21] ), .QN(n2967) );
  AO221X1 U4129 ( .IN1(n1697), .IN2(\read_value_mux[17][12] ), .IN3(
        \read_value_mux[17][21] ), .IN4(n1721), .IN5(n2967), .Q(n2973) );
  MUX21X1 U4130 ( .IN1(n1675), .IN2(search_data[5]), .S(
        \read_value_mux[17][5] ), .Q(n2971) );
  MUX21X1 U4131 ( .IN1(n1725), .IN2(search_data[23]), .S(
        \read_value_mux[17][23] ), .Q(n2970) );
  MUX21X1 U4132 ( .IN1(n1693), .IN2(search_data[11]), .S(
        \read_value_mux[17][11] ), .Q(n2969) );
  MUX21X1 U4133 ( .IN1(n1663), .IN2(search_data[1]), .S(
        \read_value_mux[17][1] ), .Q(n2968) );
  NAND4X0 U4134 ( .IN1(n2971), .IN2(n2970), .IN3(n2969), .IN4(n2968), .QN(
        n2972) );
  NOR4X0 U4135 ( .IN1(n2975), .IN2(n2974), .IN3(n2973), .IN4(n2972), .QN(n3007) );
  AOI22X1 U4136 ( .IN1(n1683), .IN2(\read_value_mux[17][7] ), .IN3(n1713), 
        .IN4(\read_value_mux[17][18] ), .QN(n2976) );
  OA221X1 U4137 ( .IN1(n1683), .IN2(\read_value_mux[17][7] ), .IN3(n1712), 
        .IN4(\read_value_mux[17][18] ), .IN5(n2976), .Q(n3006) );
  MUX21X1 U4138 ( .IN1(search_data[2]), .IN2(n1666), .S(
        \read_value_mux[17][2] ), .Q(n2983) );
  MUX21X1 U4139 ( .IN1(search_data[31]), .IN2(n1740), .S(
        \read_value_mux[17][31] ), .Q(n2982) );
  MUX21X1 U4140 ( .IN1(n1701), .IN2(search_data[14]), .S(
        \read_value_mux[17][14] ), .Q(n2980) );
  MUX21X1 U4141 ( .IN1(n1672), .IN2(search_data[4]), .S(
        \read_value_mux[17][4] ), .Q(n2979) );
  MUX21X1 U4142 ( .IN1(n1728), .IN2(search_data[26]), .S(
        \read_value_mux[17][26] ), .Q(n2978) );
  MUX21X1 U4143 ( .IN1(n1708), .IN2(search_data[16]), .S(
        \read_value_mux[17][16] ), .Q(n2977) );
  NAND4X0 U4144 ( .IN1(n2980), .IN2(n2979), .IN3(n2978), .IN4(n2977), .QN(
        n2981) );
  NOR4X0 U4145 ( .IN1(n2983), .IN2(n2982), .IN3(n1611), .IN4(n2981), .QN(n3005) );
  MUX21X1 U4146 ( .IN1(n1698), .IN2(search_data[13]), .S(
        \read_value_mux[17][13] ), .Q(n2987) );
  MUX21X1 U4147 ( .IN1(n1705), .IN2(n1704), .S(\read_value_mux[17][15] ), .Q(
        n2986) );
  MUX21X1 U4148 ( .IN1(n1717), .IN2(search_data[19]), .S(
        \read_value_mux[17][19] ), .Q(n2985) );
  MUX21X1 U4149 ( .IN1(n1718), .IN2(search_data[20]), .S(
        \read_value_mux[17][20] ), .Q(n2984) );
  NAND4X0 U4150 ( .IN1(n2987), .IN2(n2986), .IN3(n2985), .IN4(n2984), .QN(
        n3003) );
  MUX21X1 U4151 ( .IN1(n1722), .IN2(search_data[22]), .S(
        \read_value_mux[17][22] ), .Q(n2991) );
  MUX21X1 U4152 ( .IN1(n1734), .IN2(search_data[29]), .S(
        \read_value_mux[17][29] ), .Q(n2990) );
  MUX21X1 U4153 ( .IN1(n1737), .IN2(search_data[30]), .S(
        \read_value_mux[17][30] ), .Q(n2989) );
  MUX21X1 U4154 ( .IN1(n1730), .IN2(search_data[27]), .S(
        \read_value_mux[17][27] ), .Q(n2988) );
  NAND4X0 U4155 ( .IN1(n2991), .IN2(n2990), .IN3(n2989), .IN4(n2988), .QN(
        n3002) );
  MUX21X1 U4156 ( .IN1(n1733), .IN2(search_data[28]), .S(
        \read_value_mux[17][28] ), .Q(n2995) );
  MUX21X1 U4157 ( .IN1(n1662), .IN2(search_data[0]), .S(
        \read_value_mux[17][0] ), .Q(n2994) );
  MUX21X1 U4158 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[17][25] ), .Q(n2993) );
  MUX21X1 U4159 ( .IN1(n1684), .IN2(search_data[8]), .S(
        \read_value_mux[17][8] ), .Q(n2992) );
  NAND4X0 U4160 ( .IN1(n2995), .IN2(n2994), .IN3(n2993), .IN4(n2992), .QN(
        n3001) );
  MUX21X1 U4161 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[17][24] ), .Q(n2999) );
  MUX21X1 U4162 ( .IN1(n1691), .IN2(search_data[10]), .S(
        \read_value_mux[17][10] ), .Q(n2998) );
  MUX21X1 U4163 ( .IN1(n1678), .IN2(search_data[6]), .S(
        \read_value_mux[17][6] ), .Q(n2997) );
  MUX21X1 U4164 ( .IN1(n1687), .IN2(search_data[9]), .S(
        \read_value_mux[17][9] ), .Q(n2996) );
  NAND4X0 U4165 ( .IN1(n2999), .IN2(n2998), .IN3(n2997), .IN4(n2996), .QN(
        n3000) );
  NOR4X0 U4166 ( .IN1(n3003), .IN2(n3002), .IN3(n3001), .IN4(n3000), .QN(n3004) );
  NAND4X0 U4167 ( .IN1(n3007), .IN2(n3006), .IN3(n3005), .IN4(n3004), .QN(
        n3113) );
  INVX0 U4168 ( .INP(n3008), .ZN(n3009) );
  OA22X1 U4169 ( .IN1(n3064), .IN2(n3010), .IN3(n3113), .IN4(n3009), .Q(n3011)
         );
  INVX0 U4170 ( .INP(n3056), .ZN(n3120) );
  INVX0 U4171 ( .INP(n3013), .ZN(n3119) );
  NOR2X0 U4172 ( .IN1(n3120), .IN2(n3119), .QN(n3055) );
  MUX21X1 U4173 ( .IN1(search_data[15]), .IN2(n1706), .S(
        \read_value_mux[8][15] ), .Q(n3022) );
  MUX21X1 U4174 ( .IN1(search_data[30]), .IN2(n1737), .S(
        \read_value_mux[8][30] ), .Q(n3021) );
  OAI22X1 U4175 ( .IN1(\read_value_mux[8][19] ), .IN2(n1716), .IN3(n1713), 
        .IN4(\read_value_mux[8][18] ), .QN(n3014) );
  AO221X1 U4176 ( .IN1(n1717), .IN2(\read_value_mux[8][19] ), .IN3(n1714), 
        .IN4(\read_value_mux[8][18] ), .IN5(n3014), .Q(n3020) );
  MUX21X1 U4177 ( .IN1(n1682), .IN2(search_data[7]), .S(\read_value_mux[8][7] ), .Q(n3018) );
  MUX21X1 U4178 ( .IN1(n1723), .IN2(search_data[22]), .S(
        \read_value_mux[8][22] ), .Q(n3017) );
  MUX21X1 U4179 ( .IN1(n1696), .IN2(search_data[12]), .S(
        \read_value_mux[8][12] ), .Q(n3016) );
  MUX21X1 U4180 ( .IN1(n1670), .IN2(search_data[3]), .S(\read_value_mux[8][3] ), .Q(n3015) );
  NAND4X0 U4181 ( .IN1(n3018), .IN2(n3017), .IN3(n3016), .IN4(n3015), .QN(
        n3019) );
  NOR4X0 U4182 ( .IN1(n3022), .IN2(n3021), .IN3(n3020), .IN4(n3019), .QN(n3054) );
  AOI22X1 U4183 ( .IN1(n1725), .IN2(\read_value_mux[8][23] ), .IN3(n1728), 
        .IN4(\read_value_mux[8][26] ), .QN(n3023) );
  OA221X1 U4184 ( .IN1(n1725), .IN2(\read_value_mux[8][23] ), .IN3(n1729), 
        .IN4(\read_value_mux[8][26] ), .IN5(n3023), .Q(n3053) );
  MUX21X1 U4185 ( .IN1(search_data[11]), .IN2(n1693), .S(
        \read_value_mux[8][11] ), .Q(n3030) );
  MUX21X1 U4186 ( .IN1(search_data[21]), .IN2(n1719), .S(
        \read_value_mux[8][21] ), .Q(n3029) );
  MUX21X1 U4187 ( .IN1(n1735), .IN2(search_data[29]), .S(
        \read_value_mux[8][29] ), .Q(n3027) );
  MUX21X1 U4188 ( .IN1(n1740), .IN2(search_data[31]), .S(
        \read_value_mux[8][31] ), .Q(n3026) );
  MUX21X1 U4189 ( .IN1(n1731), .IN2(search_data[27]), .S(
        \read_value_mux[8][27] ), .Q(n3025) );
  MUX21X1 U4190 ( .IN1(n1679), .IN2(search_data[6]), .S(\read_value_mux[8][6] ), .Q(n3024) );
  NAND4X0 U4191 ( .IN1(n3027), .IN2(n3026), .IN3(n3025), .IN4(n3024), .QN(
        n3028) );
  NOR4X0 U4192 ( .IN1(n3030), .IN2(n3029), .IN3(n1611), .IN4(n3028), .QN(n3052) );
  MUX21X1 U4193 ( .IN1(n1663), .IN2(search_data[1]), .S(\read_value_mux[8][1] ), .Q(n3034) );
  MUX21X1 U4194 ( .IN1(n1667), .IN2(search_data[2]), .S(\read_value_mux[8][2] ), .Q(n3033) );
  MUX21X1 U4195 ( .IN1(n1660), .IN2(search_data[0]), .S(\read_value_mux[8][0] ), .Q(n3031) );
  NAND4X0 U4196 ( .IN1(n3034), .IN2(n3033), .IN3(n3032), .IN4(n3031), .QN(
        n3050) );
  MUX21X1 U4197 ( .IN1(n1726), .IN2(search_data[24]), .S(
        \read_value_mux[8][24] ), .Q(n3038) );
  MUX21X1 U4198 ( .IN1(n1673), .IN2(search_data[4]), .S(\read_value_mux[8][4] ), .Q(n3037) );
  MUX21X1 U4199 ( .IN1(n1688), .IN2(search_data[9]), .S(\read_value_mux[8][9] ), .Q(n3036) );
  MUX21X1 U4200 ( .IN1(n1702), .IN2(search_data[14]), .S(
        \read_value_mux[8][14] ), .Q(n3035) );
  NAND4X0 U4201 ( .IN1(n3038), .IN2(n3037), .IN3(n3036), .IN4(n3035), .QN(
        n3049) );
  MUX21X1 U4202 ( .IN1(n1708), .IN2(search_data[16]), .S(
        \read_value_mux[8][16] ), .Q(n3042) );
  MUX21X1 U4203 ( .IN1(n1727), .IN2(search_data[25]), .S(
        \read_value_mux[8][25] ), .Q(n3041) );
  MUX21X1 U4204 ( .IN1(n1692), .IN2(n1690), .S(\read_value_mux[8][10] ), .Q(
        n3040) );
  MUX21X1 U4205 ( .IN1(n1699), .IN2(search_data[13]), .S(
        \read_value_mux[8][13] ), .Q(n3039) );
  NAND4X0 U4206 ( .IN1(n3042), .IN2(n3041), .IN3(n3040), .IN4(n3039), .QN(
        n3048) );
  MUX21X1 U4207 ( .IN1(n1718), .IN2(search_data[20]), .S(
        \read_value_mux[8][20] ), .Q(n3046) );
  MUX21X1 U4208 ( .IN1(n1710), .IN2(search_data[17]), .S(
        \read_value_mux[8][17] ), .Q(n3045) );
  MUX21X1 U4209 ( .IN1(n1685), .IN2(search_data[8]), .S(\read_value_mux[8][8] ), .Q(n3044) );
  MUX21X1 U4210 ( .IN1(n1676), .IN2(search_data[5]), .S(\read_value_mux[8][5] ), .Q(n3043) );
  NAND4X0 U4211 ( .IN1(n3046), .IN2(n3045), .IN3(n3044), .IN4(n3043), .QN(
        n3047) );
  NOR4X0 U4212 ( .IN1(n3050), .IN2(n3049), .IN3(n3048), .IN4(n3047), .QN(n3051) );
  NAND4X0 U4213 ( .IN1(n3054), .IN2(n3053), .IN3(n3052), .IN4(n3051), .QN(
        n3095) );
  INVX0 U4214 ( .INP(n3057), .ZN(n3059) );
  NOR2X0 U4215 ( .IN1(n3059), .IN2(n3058), .QN(n3103) );
  INVX0 U4216 ( .INP(n3103), .ZN(n3100) );
  INVX0 U4217 ( .INP(n3060), .ZN(n3062) );
  NOR2X0 U4218 ( .IN1(n3062), .IN2(n3061), .QN(n3102) );
  NOR2X0 U4219 ( .IN1(n3064), .IN2(n3063), .QN(n3104) );
  INVX0 U4220 ( .INP(n3065), .ZN(n3066) );
  INVX0 U4221 ( .INP(n3068), .ZN(n3069) );
  INVX0 U4222 ( .INP(n3107), .ZN(n3086) );
  INVX0 U4223 ( .INP(n3071), .ZN(n3073) );
  NOR2X0 U4224 ( .IN1(n3073), .IN2(n3072), .QN(n3112) );
  INVX0 U4225 ( .INP(n3077), .ZN(n3078) );
  INVX0 U4226 ( .INP(n3080), .ZN(n3110) );
  AO221X1 U4227 ( .IN1(n3112), .IN2(n1612), .IN3(n3112), .IN4(n3109), .IN5(
        n3081), .Q(n3085) );
  INVX0 U4228 ( .INP(n3082), .ZN(n3084) );
  NOR2X0 U4229 ( .IN1(n3084), .IN2(n3083), .QN(n3115) );
  OA221X1 U4230 ( .IN1(n3108), .IN2(n3086), .IN3(n3108), .IN4(n3085), .IN5(
        n3115), .Q(n3092) );
  INVX0 U4231 ( .INP(n3087), .ZN(n3114) );
  INVX0 U4232 ( .INP(n3088), .ZN(n3090) );
  NOR2X0 U4233 ( .IN1(n3090), .IN2(n3089), .QN(n3125) );
  OA21X1 U4234 ( .IN1(n3092), .IN2(n3091), .IN3(n3125), .Q(n3097) );
  INVX0 U4235 ( .INP(n3093), .ZN(n3122) );
  AO221X1 U4236 ( .IN1(n3104), .IN2(n3097), .IN3(n3104), .IN4(n3096), .IN5(
        n3106), .Q(n3099) );
  NOR2X0 U4237 ( .IN1(n3119), .IN2(n3117), .QN(n3098) );
  OA221X1 U4238 ( .IN1(n3100), .IN2(n3102), .IN3(n3100), .IN4(n3099), .IN5(
        n3098), .Q(n3101) );
  INVX0 U4239 ( .INP(n3104), .ZN(n3105) );
  NOR2X0 U4240 ( .IN1(n3106), .IN2(n3105), .QN(n3124) );
  NOR2X0 U4241 ( .IN1(n3108), .IN2(n3107), .QN(n3127) );
  NAND3X0 U4242 ( .IN1(n3115), .IN2(n3114), .IN3(n3113), .QN(n3126) );
  AO221X1 U4243 ( .IN1(n3127), .IN2(n3130), .IN3(n3127), .IN4(n3129), .IN5(
        n3126), .Q(n3116) );
  NAND4X0 U4244 ( .IN1(n3125), .IN2(n3123), .IN3(n3122), .IN4(n3116), .QN(
        n3121) );
  NOR4X0 U4245 ( .IN1(n3120), .IN2(n3119), .IN3(n3118), .IN4(n3117), .QN(n3132) );
  OA221X1 U4246 ( .IN1(n3137), .IN2(n3124), .IN3(n3137), .IN4(n3121), .IN5(
        n3132), .Q(search_index[2]) );
  NAND4X0 U4247 ( .IN1(n3125), .IN2(n3124), .IN3(n3123), .IN4(n3122), .QN(
        n3139) );
  INVX0 U4248 ( .INP(n3126), .ZN(n3128) );
  INVX0 U4249 ( .INP(n3135), .ZN(n3133) );
  INVX0 U4250 ( .INP(n3129), .ZN(n3131) );
  INVX0 U4251 ( .INP(n3132), .ZN(n3136) );
  NOR2X0 U4252 ( .IN1(n3136), .IN2(n3137), .QN(n3138) );
  OA221X1 U4253 ( .IN1(n3139), .IN2(n3133), .IN3(n3139), .IN4(n3134), .IN5(
        n3138), .Q(search_index[3]) );
  NOR2X0 U4254 ( .IN1(n3135), .IN2(n3134), .QN(n3140) );
  NOR4X0 U4255 ( .IN1(n3140), .IN2(n3137), .IN3(n3136), .IN4(n3139), .QN(
        search_index[4]) );
  AO22X1 U4256 ( .IN1(\read_value_mux[0][0] ), .IN2(n1617), .IN3(write_data[0]), .IN4(n3141), .Q(\words[0]/data_i[0] ) );
  AO22X1 U4257 ( .IN1(\read_value_mux[0][10] ), .IN2(n1617), .IN3(n3141), 
        .IN4(write_data[10]), .Q(\words[0]/data_i[10] ) );
  AO22X1 U4258 ( .IN1(\read_value_mux[0][11] ), .IN2(n1617), .IN3(n3141), 
        .IN4(write_data[11]), .Q(\words[0]/data_i[11] ) );
  AO22X1 U4259 ( .IN1(\read_value_mux[0][12] ), .IN2(n1617), .IN3(n3141), 
        .IN4(write_data[12]), .Q(\words[0]/data_i[12] ) );
  AO22X1 U4260 ( .IN1(\read_value_mux[0][13] ), .IN2(n1617), .IN3(n3141), 
        .IN4(write_data[13]), .Q(\words[0]/data_i[13] ) );
  AO22X1 U4261 ( .IN1(\read_value_mux[0][14] ), .IN2(n1617), .IN3(n3141), 
        .IN4(write_data[14]), .Q(\words[0]/data_i[14] ) );
  AO22X1 U4262 ( .IN1(\read_value_mux[0][15] ), .IN2(n1617), .IN3(n3141), 
        .IN4(write_data[15]), .Q(\words[0]/data_i[15] ) );
  AO22X1 U4263 ( .IN1(\read_value_mux[0][16] ), .IN2(n1617), .IN3(n3141), 
        .IN4(write_data[16]), .Q(\words[0]/data_i[16] ) );
  AO22X1 U4264 ( .IN1(\read_value_mux[0][17] ), .IN2(n1617), .IN3(n3141), 
        .IN4(write_data[17]), .Q(\words[0]/data_i[17] ) );
  AO22X1 U4265 ( .IN1(\read_value_mux[0][18] ), .IN2(n1617), .IN3(n3141), 
        .IN4(write_data[18]), .Q(\words[0]/data_i[18] ) );
  AO22X1 U4266 ( .IN1(\read_value_mux[0][19] ), .IN2(n1617), .IN3(n3141), 
        .IN4(write_data[19]), .Q(\words[0]/data_i[19] ) );
  AO22X1 U4267 ( .IN1(\read_value_mux[0][1] ), .IN2(n1617), .IN3(n3141), .IN4(
        write_data[1]), .Q(\words[0]/data_i[1] ) );
  AO22X1 U4268 ( .IN1(\read_value_mux[0][20] ), .IN2(n1617), .IN3(n3141), 
        .IN4(write_data[20]), .Q(\words[0]/data_i[20] ) );
  AO22X1 U4269 ( .IN1(\read_value_mux[0][21] ), .IN2(n1617), .IN3(n3141), 
        .IN4(write_data[21]), .Q(\words[0]/data_i[21] ) );
  AO22X1 U4270 ( .IN1(\read_value_mux[0][22] ), .IN2(n1617), .IN3(n3141), 
        .IN4(write_data[22]), .Q(\words[0]/data_i[22] ) );
  AO22X1 U4271 ( .IN1(\read_value_mux[0][23] ), .IN2(n1617), .IN3(n3141), 
        .IN4(write_data[23]), .Q(\words[0]/data_i[23] ) );
  AO22X1 U4272 ( .IN1(\read_value_mux[0][24] ), .IN2(n1617), .IN3(n3141), 
        .IN4(write_data[24]), .Q(\words[0]/data_i[24] ) );
  AO22X1 U4273 ( .IN1(\read_value_mux[0][25] ), .IN2(n1617), .IN3(n3141), 
        .IN4(write_data[25]), .Q(\words[0]/data_i[25] ) );
  AO22X1 U4274 ( .IN1(\read_value_mux[0][26] ), .IN2(n1617), .IN3(n3141), 
        .IN4(write_data[26]), .Q(\words[0]/data_i[26] ) );
  AO22X1 U4275 ( .IN1(\read_value_mux[0][27] ), .IN2(n1617), .IN3(n3141), 
        .IN4(write_data[27]), .Q(\words[0]/data_i[27] ) );
  AO22X1 U4276 ( .IN1(\read_value_mux[0][28] ), .IN2(n1617), .IN3(n3141), 
        .IN4(write_data[28]), .Q(\words[0]/data_i[28] ) );
  AO22X1 U4277 ( .IN1(\read_value_mux[0][29] ), .IN2(n1617), .IN3(n3141), 
        .IN4(write_data[29]), .Q(\words[0]/data_i[29] ) );
  AO22X1 U4278 ( .IN1(\read_value_mux[0][2] ), .IN2(n1617), .IN3(n3141), .IN4(
        write_data[2]), .Q(\words[0]/data_i[2] ) );
  AO22X1 U4279 ( .IN1(\read_value_mux[0][30] ), .IN2(n1617), .IN3(n3141), 
        .IN4(write_data[30]), .Q(\words[0]/data_i[30] ) );
  AO22X1 U4280 ( .IN1(\read_value_mux[0][31] ), .IN2(n1617), .IN3(n3141), 
        .IN4(write_data[31]), .Q(\words[0]/data_i[31] ) );
  AO22X1 U4281 ( .IN1(\read_value_mux[0][3] ), .IN2(n1617), .IN3(n3141), .IN4(
        write_data[3]), .Q(\words[0]/data_i[3] ) );
  AO22X1 U4282 ( .IN1(\read_value_mux[0][4] ), .IN2(n1617), .IN3(n3141), .IN4(
        write_data[4]), .Q(\words[0]/data_i[4] ) );
  AO22X1 U4283 ( .IN1(\read_value_mux[0][5] ), .IN2(n1617), .IN3(n3141), .IN4(
        write_data[5]), .Q(\words[0]/data_i[5] ) );
  AO22X1 U4284 ( .IN1(\read_value_mux[0][6] ), .IN2(n1617), .IN3(n3141), .IN4(
        write_data[6]), .Q(\words[0]/data_i[6] ) );
  AO22X1 U4285 ( .IN1(\read_value_mux[0][7] ), .IN2(n1617), .IN3(n3141), .IN4(
        write_data[7]), .Q(\words[0]/data_i[7] ) );
  AO22X1 U4286 ( .IN1(\read_value_mux[0][8] ), .IN2(n1617), .IN3(n3141), .IN4(
        write_data[8]), .Q(\words[0]/data_i[8] ) );
  AO22X1 U4287 ( .IN1(\read_value_mux[0][9] ), .IN2(n1617), .IN3(n3141), .IN4(
        write_data[9]), .Q(\words[0]/data_i[9] ) );
  AO21X1 U4288 ( .IN1(\words[0]/valid_o ), .IN2(n1743), .IN3(n3141), .Q(
        \words[0]/valid_i ) );
  AO22X1 U4289 ( .IN1(\read_value_mux[10][0] ), .IN2(n1614), .IN3(
        write_data[0]), .IN4(n3142), .Q(\words[10]/data_i[0] ) );
  AO22X1 U4290 ( .IN1(\read_value_mux[10][10] ), .IN2(n1614), .IN3(
        write_data[10]), .IN4(n3142), .Q(\words[10]/data_i[10] ) );
  AO22X1 U4291 ( .IN1(\read_value_mux[10][11] ), .IN2(n1614), .IN3(
        write_data[11]), .IN4(n3142), .Q(\words[10]/data_i[11] ) );
  AO22X1 U4292 ( .IN1(\read_value_mux[10][12] ), .IN2(n1614), .IN3(
        write_data[12]), .IN4(n3142), .Q(\words[10]/data_i[12] ) );
  AO22X1 U4293 ( .IN1(\read_value_mux[10][13] ), .IN2(n1614), .IN3(
        write_data[13]), .IN4(n3142), .Q(\words[10]/data_i[13] ) );
  AO22X1 U4294 ( .IN1(\read_value_mux[10][14] ), .IN2(n1614), .IN3(
        write_data[14]), .IN4(n3142), .Q(\words[10]/data_i[14] ) );
  AO22X1 U4295 ( .IN1(\read_value_mux[10][15] ), .IN2(n1614), .IN3(
        write_data[15]), .IN4(n3142), .Q(\words[10]/data_i[15] ) );
  AO22X1 U4296 ( .IN1(\read_value_mux[10][16] ), .IN2(n1614), .IN3(
        write_data[16]), .IN4(n3142), .Q(\words[10]/data_i[16] ) );
  AO22X1 U4297 ( .IN1(\read_value_mux[10][17] ), .IN2(n1614), .IN3(
        write_data[17]), .IN4(n3142), .Q(\words[10]/data_i[17] ) );
  AO22X1 U4298 ( .IN1(\read_value_mux[10][18] ), .IN2(n1614), .IN3(
        write_data[18]), .IN4(n3142), .Q(\words[10]/data_i[18] ) );
  AO22X1 U4299 ( .IN1(\read_value_mux[10][19] ), .IN2(n1614), .IN3(
        write_data[19]), .IN4(n3142), .Q(\words[10]/data_i[19] ) );
  AO22X1 U4300 ( .IN1(\read_value_mux[10][1] ), .IN2(n1614), .IN3(
        write_data[1]), .IN4(n3142), .Q(\words[10]/data_i[1] ) );
  AO22X1 U4301 ( .IN1(\read_value_mux[10][20] ), .IN2(n1614), .IN3(
        write_data[20]), .IN4(n3142), .Q(\words[10]/data_i[20] ) );
  AO22X1 U4302 ( .IN1(\read_value_mux[10][21] ), .IN2(n1614), .IN3(
        write_data[21]), .IN4(n3142), .Q(\words[10]/data_i[21] ) );
  AO22X1 U4303 ( .IN1(\read_value_mux[10][22] ), .IN2(n1614), .IN3(
        write_data[22]), .IN4(n3142), .Q(\words[10]/data_i[22] ) );
  AO22X1 U4304 ( .IN1(\read_value_mux[10][23] ), .IN2(n1614), .IN3(
        write_data[23]), .IN4(n3142), .Q(\words[10]/data_i[23] ) );
  AO22X1 U4305 ( .IN1(\read_value_mux[10][24] ), .IN2(n1614), .IN3(
        write_data[24]), .IN4(n3142), .Q(\words[10]/data_i[24] ) );
  AO22X1 U4306 ( .IN1(\read_value_mux[10][25] ), .IN2(n1614), .IN3(
        write_data[25]), .IN4(n3142), .Q(\words[10]/data_i[25] ) );
  AO22X1 U4307 ( .IN1(\read_value_mux[10][26] ), .IN2(n1614), .IN3(
        write_data[26]), .IN4(n3142), .Q(\words[10]/data_i[26] ) );
  AO22X1 U4308 ( .IN1(\read_value_mux[10][27] ), .IN2(n1614), .IN3(
        write_data[27]), .IN4(n3142), .Q(\words[10]/data_i[27] ) );
  AO22X1 U4309 ( .IN1(\read_value_mux[10][28] ), .IN2(n1614), .IN3(
        write_data[28]), .IN4(n3142), .Q(\words[10]/data_i[28] ) );
  AO22X1 U4310 ( .IN1(\read_value_mux[10][29] ), .IN2(n1614), .IN3(
        write_data[29]), .IN4(n3142), .Q(\words[10]/data_i[29] ) );
  AO22X1 U4311 ( .IN1(\read_value_mux[10][2] ), .IN2(n1614), .IN3(
        write_data[2]), .IN4(n3142), .Q(\words[10]/data_i[2] ) );
  AO22X1 U4312 ( .IN1(\read_value_mux[10][30] ), .IN2(n1614), .IN3(
        write_data[30]), .IN4(n3142), .Q(\words[10]/data_i[30] ) );
  AO22X1 U4313 ( .IN1(\read_value_mux[10][31] ), .IN2(n1614), .IN3(
        write_data[31]), .IN4(n3142), .Q(\words[10]/data_i[31] ) );
  AO22X1 U4314 ( .IN1(\read_value_mux[10][3] ), .IN2(n1614), .IN3(
        write_data[3]), .IN4(n3142), .Q(\words[10]/data_i[3] ) );
  AO22X1 U4315 ( .IN1(\read_value_mux[10][4] ), .IN2(n1614), .IN3(
        write_data[4]), .IN4(n3142), .Q(\words[10]/data_i[4] ) );
  AO22X1 U4316 ( .IN1(\read_value_mux[10][5] ), .IN2(n1614), .IN3(
        write_data[5]), .IN4(n3142), .Q(\words[10]/data_i[5] ) );
  AO22X1 U4317 ( .IN1(\read_value_mux[10][6] ), .IN2(n1614), .IN3(
        write_data[6]), .IN4(n3142), .Q(\words[10]/data_i[6] ) );
  AO22X1 U4318 ( .IN1(\read_value_mux[10][7] ), .IN2(n1614), .IN3(
        write_data[7]), .IN4(n3142), .Q(\words[10]/data_i[7] ) );
  AO22X1 U4319 ( .IN1(\read_value_mux[10][8] ), .IN2(n1614), .IN3(
        write_data[8]), .IN4(n3142), .Q(\words[10]/data_i[8] ) );
  AO22X1 U4320 ( .IN1(\read_value_mux[10][9] ), .IN2(n1614), .IN3(
        write_data[9]), .IN4(n3142), .Q(\words[10]/data_i[9] ) );
  AO21X1 U4321 ( .IN1(\words[10]/valid_o ), .IN2(n1743), .IN3(n3142), .Q(
        \words[10]/valid_i ) );
  AO22X1 U4322 ( .IN1(\read_value_mux[11][0] ), .IN2(n1623), .IN3(
        write_data[0]), .IN4(n3143), .Q(\words[11]/data_i[0] ) );
  AO22X1 U4323 ( .IN1(\read_value_mux[11][10] ), .IN2(n1623), .IN3(
        write_data[10]), .IN4(n3143), .Q(\words[11]/data_i[10] ) );
  AO22X1 U4324 ( .IN1(\read_value_mux[11][11] ), .IN2(n1623), .IN3(
        write_data[11]), .IN4(n3143), .Q(\words[11]/data_i[11] ) );
  AO22X1 U4325 ( .IN1(\read_value_mux[11][12] ), .IN2(n1623), .IN3(
        write_data[12]), .IN4(n3143), .Q(\words[11]/data_i[12] ) );
  AO22X1 U4326 ( .IN1(\read_value_mux[11][13] ), .IN2(n1623), .IN3(
        write_data[13]), .IN4(n3143), .Q(\words[11]/data_i[13] ) );
  AO22X1 U4327 ( .IN1(\read_value_mux[11][14] ), .IN2(n1623), .IN3(
        write_data[14]), .IN4(n3143), .Q(\words[11]/data_i[14] ) );
  AO22X1 U4328 ( .IN1(\read_value_mux[11][15] ), .IN2(n1623), .IN3(
        write_data[15]), .IN4(n3143), .Q(\words[11]/data_i[15] ) );
  AO22X1 U4329 ( .IN1(\read_value_mux[11][16] ), .IN2(n1623), .IN3(
        write_data[16]), .IN4(n3143), .Q(\words[11]/data_i[16] ) );
  AO22X1 U4330 ( .IN1(\read_value_mux[11][17] ), .IN2(n1623), .IN3(
        write_data[17]), .IN4(n3143), .Q(\words[11]/data_i[17] ) );
  AO22X1 U4331 ( .IN1(\read_value_mux[11][18] ), .IN2(n1623), .IN3(
        write_data[18]), .IN4(n3143), .Q(\words[11]/data_i[18] ) );
  AO22X1 U4332 ( .IN1(\read_value_mux[11][19] ), .IN2(n1623), .IN3(
        write_data[19]), .IN4(n3143), .Q(\words[11]/data_i[19] ) );
  AO22X1 U4333 ( .IN1(\read_value_mux[11][1] ), .IN2(n1623), .IN3(
        write_data[1]), .IN4(n3143), .Q(\words[11]/data_i[1] ) );
  AO22X1 U4334 ( .IN1(\read_value_mux[11][20] ), .IN2(n1623), .IN3(
        write_data[20]), .IN4(n3143), .Q(\words[11]/data_i[20] ) );
  AO22X1 U4335 ( .IN1(\read_value_mux[11][21] ), .IN2(n1623), .IN3(
        write_data[21]), .IN4(n3143), .Q(\words[11]/data_i[21] ) );
  AO22X1 U4336 ( .IN1(\read_value_mux[11][22] ), .IN2(n1623), .IN3(
        write_data[22]), .IN4(n3143), .Q(\words[11]/data_i[22] ) );
  AO22X1 U4337 ( .IN1(\read_value_mux[11][23] ), .IN2(n1623), .IN3(
        write_data[23]), .IN4(n3143), .Q(\words[11]/data_i[23] ) );
  AO22X1 U4338 ( .IN1(\read_value_mux[11][24] ), .IN2(n1623), .IN3(
        write_data[24]), .IN4(n3143), .Q(\words[11]/data_i[24] ) );
  AO22X1 U4339 ( .IN1(\read_value_mux[11][25] ), .IN2(n1623), .IN3(
        write_data[25]), .IN4(n3143), .Q(\words[11]/data_i[25] ) );
  AO22X1 U4340 ( .IN1(\read_value_mux[11][26] ), .IN2(n1623), .IN3(
        write_data[26]), .IN4(n3143), .Q(\words[11]/data_i[26] ) );
  AO22X1 U4341 ( .IN1(\read_value_mux[11][27] ), .IN2(n1623), .IN3(
        write_data[27]), .IN4(n3143), .Q(\words[11]/data_i[27] ) );
  AO22X1 U4342 ( .IN1(\read_value_mux[11][28] ), .IN2(n1623), .IN3(
        write_data[28]), .IN4(n3143), .Q(\words[11]/data_i[28] ) );
  AO22X1 U4343 ( .IN1(\read_value_mux[11][29] ), .IN2(n1623), .IN3(
        write_data[29]), .IN4(n3143), .Q(\words[11]/data_i[29] ) );
  AO22X1 U4344 ( .IN1(\read_value_mux[11][2] ), .IN2(n1623), .IN3(
        write_data[2]), .IN4(n3143), .Q(\words[11]/data_i[2] ) );
  AO22X1 U4345 ( .IN1(\read_value_mux[11][30] ), .IN2(n1623), .IN3(
        write_data[30]), .IN4(n3143), .Q(\words[11]/data_i[30] ) );
  AO22X1 U4346 ( .IN1(\read_value_mux[11][31] ), .IN2(n1623), .IN3(
        write_data[31]), .IN4(n3143), .Q(\words[11]/data_i[31] ) );
  AO22X1 U4347 ( .IN1(\read_value_mux[11][3] ), .IN2(n1623), .IN3(
        write_data[3]), .IN4(n3143), .Q(\words[11]/data_i[3] ) );
  AO22X1 U4348 ( .IN1(\read_value_mux[11][4] ), .IN2(n1623), .IN3(
        write_data[4]), .IN4(n3143), .Q(\words[11]/data_i[4] ) );
  AO22X1 U4349 ( .IN1(\read_value_mux[11][5] ), .IN2(n1623), .IN3(
        write_data[5]), .IN4(n3143), .Q(\words[11]/data_i[5] ) );
  AO22X1 U4350 ( .IN1(\read_value_mux[11][6] ), .IN2(n1623), .IN3(
        write_data[6]), .IN4(n3143), .Q(\words[11]/data_i[6] ) );
  AO22X1 U4351 ( .IN1(\read_value_mux[11][7] ), .IN2(n1623), .IN3(
        write_data[7]), .IN4(n3143), .Q(\words[11]/data_i[7] ) );
  AO22X1 U4352 ( .IN1(\read_value_mux[11][8] ), .IN2(n1623), .IN3(
        write_data[8]), .IN4(n3143), .Q(\words[11]/data_i[8] ) );
  AO22X1 U4353 ( .IN1(\read_value_mux[11][9] ), .IN2(n1623), .IN3(
        write_data[9]), .IN4(n3143), .Q(\words[11]/data_i[9] ) );
  AO21X1 U4354 ( .IN1(\words[11]/valid_o ), .IN2(n1743), .IN3(n3143), .Q(
        \words[11]/valid_i ) );
  AO22X1 U4355 ( .IN1(\read_value_mux[12][0] ), .IN2(n1618), .IN3(
        write_data[0]), .IN4(n3144), .Q(\words[12]/data_i[0] ) );
  AO22X1 U4356 ( .IN1(\read_value_mux[12][10] ), .IN2(n1618), .IN3(
        write_data[10]), .IN4(n3144), .Q(\words[12]/data_i[10] ) );
  AO22X1 U4357 ( .IN1(\read_value_mux[12][11] ), .IN2(n1618), .IN3(
        write_data[11]), .IN4(n3144), .Q(\words[12]/data_i[11] ) );
  AO22X1 U4358 ( .IN1(\read_value_mux[12][12] ), .IN2(n1618), .IN3(
        write_data[12]), .IN4(n3144), .Q(\words[12]/data_i[12] ) );
  AO22X1 U4359 ( .IN1(\read_value_mux[12][13] ), .IN2(n1618), .IN3(
        write_data[13]), .IN4(n3144), .Q(\words[12]/data_i[13] ) );
  AO22X1 U4360 ( .IN1(\read_value_mux[12][14] ), .IN2(n1618), .IN3(
        write_data[14]), .IN4(n3144), .Q(\words[12]/data_i[14] ) );
  AO22X1 U4361 ( .IN1(\read_value_mux[12][15] ), .IN2(n1618), .IN3(
        write_data[15]), .IN4(n3144), .Q(\words[12]/data_i[15] ) );
  AO22X1 U4362 ( .IN1(\read_value_mux[12][16] ), .IN2(n1618), .IN3(
        write_data[16]), .IN4(n3144), .Q(\words[12]/data_i[16] ) );
  AO22X1 U4363 ( .IN1(\read_value_mux[12][17] ), .IN2(n1618), .IN3(
        write_data[17]), .IN4(n3144), .Q(\words[12]/data_i[17] ) );
  AO22X1 U4364 ( .IN1(\read_value_mux[12][18] ), .IN2(n1618), .IN3(
        write_data[18]), .IN4(n3144), .Q(\words[12]/data_i[18] ) );
  AO22X1 U4365 ( .IN1(\read_value_mux[12][19] ), .IN2(n1618), .IN3(
        write_data[19]), .IN4(n3144), .Q(\words[12]/data_i[19] ) );
  AO22X1 U4366 ( .IN1(\read_value_mux[12][1] ), .IN2(n1618), .IN3(
        write_data[1]), .IN4(n3144), .Q(\words[12]/data_i[1] ) );
  AO22X1 U4367 ( .IN1(\read_value_mux[12][20] ), .IN2(n1618), .IN3(
        write_data[20]), .IN4(n3144), .Q(\words[12]/data_i[20] ) );
  AO22X1 U4368 ( .IN1(\read_value_mux[12][21] ), .IN2(n1618), .IN3(
        write_data[21]), .IN4(n3144), .Q(\words[12]/data_i[21] ) );
  AO22X1 U4369 ( .IN1(\read_value_mux[12][22] ), .IN2(n1618), .IN3(
        write_data[22]), .IN4(n3144), .Q(\words[12]/data_i[22] ) );
  AO22X1 U4370 ( .IN1(\read_value_mux[12][23] ), .IN2(n1618), .IN3(
        write_data[23]), .IN4(n3144), .Q(\words[12]/data_i[23] ) );
  AO22X1 U4371 ( .IN1(\read_value_mux[12][24] ), .IN2(n1618), .IN3(
        write_data[24]), .IN4(n3144), .Q(\words[12]/data_i[24] ) );
  AO22X1 U4372 ( .IN1(\read_value_mux[12][25] ), .IN2(n1618), .IN3(
        write_data[25]), .IN4(n3144), .Q(\words[12]/data_i[25] ) );
  AO22X1 U4373 ( .IN1(\read_value_mux[12][26] ), .IN2(n1618), .IN3(
        write_data[26]), .IN4(n3144), .Q(\words[12]/data_i[26] ) );
  AO22X1 U4374 ( .IN1(\read_value_mux[12][27] ), .IN2(n1618), .IN3(
        write_data[27]), .IN4(n3144), .Q(\words[12]/data_i[27] ) );
  AO22X1 U4375 ( .IN1(\read_value_mux[12][28] ), .IN2(n1618), .IN3(
        write_data[28]), .IN4(n3144), .Q(\words[12]/data_i[28] ) );
  AO22X1 U4376 ( .IN1(\read_value_mux[12][29] ), .IN2(n1618), .IN3(
        write_data[29]), .IN4(n3144), .Q(\words[12]/data_i[29] ) );
  AO22X1 U4377 ( .IN1(\read_value_mux[12][2] ), .IN2(n1618), .IN3(
        write_data[2]), .IN4(n3144), .Q(\words[12]/data_i[2] ) );
  AO22X1 U4378 ( .IN1(\read_value_mux[12][30] ), .IN2(n1618), .IN3(
        write_data[30]), .IN4(n3144), .Q(\words[12]/data_i[30] ) );
  AO22X1 U4379 ( .IN1(\read_value_mux[12][31] ), .IN2(n1618), .IN3(
        write_data[31]), .IN4(n3144), .Q(\words[12]/data_i[31] ) );
  AO22X1 U4380 ( .IN1(\read_value_mux[12][3] ), .IN2(n1618), .IN3(
        write_data[3]), .IN4(n3144), .Q(\words[12]/data_i[3] ) );
  AO22X1 U4381 ( .IN1(\read_value_mux[12][4] ), .IN2(n1618), .IN3(
        write_data[4]), .IN4(n3144), .Q(\words[12]/data_i[4] ) );
  AO22X1 U4382 ( .IN1(\read_value_mux[12][5] ), .IN2(n1618), .IN3(
        write_data[5]), .IN4(n3144), .Q(\words[12]/data_i[5] ) );
  AO22X1 U4383 ( .IN1(\read_value_mux[12][6] ), .IN2(n1618), .IN3(
        write_data[6]), .IN4(n3144), .Q(\words[12]/data_i[6] ) );
  AO22X1 U4384 ( .IN1(\read_value_mux[12][7] ), .IN2(n1618), .IN3(
        write_data[7]), .IN4(n3144), .Q(\words[12]/data_i[7] ) );
  AO22X1 U4385 ( .IN1(\read_value_mux[12][8] ), .IN2(n1618), .IN3(
        write_data[8]), .IN4(n3144), .Q(\words[12]/data_i[8] ) );
  AO22X1 U4386 ( .IN1(\read_value_mux[12][9] ), .IN2(n1618), .IN3(
        write_data[9]), .IN4(n3144), .Q(\words[12]/data_i[9] ) );
  AO21X1 U4387 ( .IN1(\words[12]/valid_o ), .IN2(n1743), .IN3(n3144), .Q(
        \words[12]/valid_i ) );
  AO22X1 U4388 ( .IN1(\read_value_mux[13][0] ), .IN2(n1619), .IN3(
        write_data[0]), .IN4(n3146), .Q(\words[13]/data_i[0] ) );
  AO22X1 U4389 ( .IN1(\read_value_mux[13][10] ), .IN2(n1619), .IN3(
        write_data[10]), .IN4(n3146), .Q(\words[13]/data_i[10] ) );
  AO22X1 U4390 ( .IN1(\read_value_mux[13][11] ), .IN2(n1619), .IN3(
        write_data[11]), .IN4(n3146), .Q(\words[13]/data_i[11] ) );
  AO22X1 U4391 ( .IN1(\read_value_mux[13][12] ), .IN2(n1619), .IN3(
        write_data[12]), .IN4(n3146), .Q(\words[13]/data_i[12] ) );
  AO22X1 U4392 ( .IN1(\read_value_mux[13][13] ), .IN2(n1619), .IN3(
        write_data[13]), .IN4(n3146), .Q(\words[13]/data_i[13] ) );
  AO22X1 U4393 ( .IN1(\read_value_mux[13][14] ), .IN2(n1619), .IN3(
        write_data[14]), .IN4(n3146), .Q(\words[13]/data_i[14] ) );
  AO22X1 U4394 ( .IN1(\read_value_mux[13][15] ), .IN2(n1619), .IN3(
        write_data[15]), .IN4(n3146), .Q(\words[13]/data_i[15] ) );
  AO22X1 U4395 ( .IN1(\read_value_mux[13][16] ), .IN2(n1619), .IN3(
        write_data[16]), .IN4(n3146), .Q(\words[13]/data_i[16] ) );
  AO22X1 U4396 ( .IN1(\read_value_mux[13][17] ), .IN2(n1619), .IN3(
        write_data[17]), .IN4(n3146), .Q(\words[13]/data_i[17] ) );
  AO22X1 U4397 ( .IN1(\read_value_mux[13][18] ), .IN2(n1619), .IN3(
        write_data[18]), .IN4(n3146), .Q(\words[13]/data_i[18] ) );
  AO22X1 U4398 ( .IN1(\read_value_mux[13][19] ), .IN2(n1619), .IN3(
        write_data[19]), .IN4(n3146), .Q(\words[13]/data_i[19] ) );
  AO22X1 U4399 ( .IN1(\read_value_mux[13][1] ), .IN2(n1619), .IN3(
        write_data[1]), .IN4(n3146), .Q(\words[13]/data_i[1] ) );
  AO22X1 U4400 ( .IN1(\read_value_mux[13][20] ), .IN2(n1619), .IN3(
        write_data[20]), .IN4(n3146), .Q(\words[13]/data_i[20] ) );
  AO22X1 U4401 ( .IN1(\read_value_mux[13][21] ), .IN2(n1619), .IN3(
        write_data[21]), .IN4(n3146), .Q(\words[13]/data_i[21] ) );
  AO22X1 U4402 ( .IN1(\read_value_mux[13][22] ), .IN2(n1619), .IN3(
        write_data[22]), .IN4(n3146), .Q(\words[13]/data_i[22] ) );
  AO22X1 U4403 ( .IN1(\read_value_mux[13][23] ), .IN2(n1619), .IN3(
        write_data[23]), .IN4(n3146), .Q(\words[13]/data_i[23] ) );
  AO22X1 U4404 ( .IN1(\read_value_mux[13][24] ), .IN2(n1619), .IN3(
        write_data[24]), .IN4(n3146), .Q(\words[13]/data_i[24] ) );
  AO22X1 U4405 ( .IN1(\read_value_mux[13][25] ), .IN2(n1619), .IN3(
        write_data[25]), .IN4(n3146), .Q(\words[13]/data_i[25] ) );
  AO22X1 U4406 ( .IN1(\read_value_mux[13][26] ), .IN2(n1619), .IN3(
        write_data[26]), .IN4(n3146), .Q(\words[13]/data_i[26] ) );
  AO22X1 U4407 ( .IN1(\read_value_mux[13][27] ), .IN2(n1619), .IN3(
        write_data[27]), .IN4(n3146), .Q(\words[13]/data_i[27] ) );
  AO22X1 U4408 ( .IN1(\read_value_mux[13][28] ), .IN2(n1619), .IN3(
        write_data[28]), .IN4(n3146), .Q(\words[13]/data_i[28] ) );
  AO22X1 U4409 ( .IN1(\read_value_mux[13][29] ), .IN2(n1619), .IN3(
        write_data[29]), .IN4(n3146), .Q(\words[13]/data_i[29] ) );
  AO22X1 U4410 ( .IN1(\read_value_mux[13][2] ), .IN2(n1619), .IN3(
        write_data[2]), .IN4(n3146), .Q(\words[13]/data_i[2] ) );
  AO22X1 U4411 ( .IN1(\read_value_mux[13][30] ), .IN2(n1619), .IN3(
        write_data[30]), .IN4(n3146), .Q(\words[13]/data_i[30] ) );
  AO22X1 U4412 ( .IN1(\read_value_mux[13][31] ), .IN2(n1619), .IN3(
        write_data[31]), .IN4(n3146), .Q(\words[13]/data_i[31] ) );
  AO22X1 U4413 ( .IN1(\read_value_mux[13][3] ), .IN2(n1619), .IN3(
        write_data[3]), .IN4(n3146), .Q(\words[13]/data_i[3] ) );
  AO22X1 U4414 ( .IN1(\read_value_mux[13][4] ), .IN2(n1619), .IN3(
        write_data[4]), .IN4(n3146), .Q(\words[13]/data_i[4] ) );
  AO22X1 U4415 ( .IN1(\read_value_mux[13][5] ), .IN2(n1619), .IN3(
        write_data[5]), .IN4(n3146), .Q(\words[13]/data_i[5] ) );
  AO22X1 U4416 ( .IN1(\read_value_mux[13][6] ), .IN2(n1619), .IN3(
        write_data[6]), .IN4(n3146), .Q(\words[13]/data_i[6] ) );
  AO22X1 U4417 ( .IN1(\read_value_mux[13][7] ), .IN2(n1619), .IN3(
        write_data[7]), .IN4(n3146), .Q(\words[13]/data_i[7] ) );
  AO22X1 U4418 ( .IN1(\read_value_mux[13][8] ), .IN2(n1619), .IN3(
        write_data[8]), .IN4(n3146), .Q(\words[13]/data_i[8] ) );
  AO22X1 U4419 ( .IN1(\read_value_mux[13][9] ), .IN2(n1619), .IN3(
        write_data[9]), .IN4(n3146), .Q(\words[13]/data_i[9] ) );
  AO21X1 U4420 ( .IN1(\words[13]/valid_o ), .IN2(n1743), .IN3(n3146), .Q(
        \words[13]/valid_i ) );
  AO22X1 U4421 ( .IN1(\read_value_mux[14][0] ), .IN2(n1624), .IN3(
        write_data[0]), .IN4(n3147), .Q(\words[14]/data_i[0] ) );
  AO22X1 U4422 ( .IN1(\read_value_mux[14][10] ), .IN2(n1624), .IN3(
        write_data[10]), .IN4(n3147), .Q(\words[14]/data_i[10] ) );
  AO22X1 U4423 ( .IN1(\read_value_mux[14][11] ), .IN2(n1624), .IN3(
        write_data[11]), .IN4(n3147), .Q(\words[14]/data_i[11] ) );
  AO22X1 U4424 ( .IN1(\read_value_mux[14][12] ), .IN2(n1624), .IN3(
        write_data[12]), .IN4(n3147), .Q(\words[14]/data_i[12] ) );
  AO22X1 U4425 ( .IN1(\read_value_mux[14][13] ), .IN2(n1624), .IN3(
        write_data[13]), .IN4(n3147), .Q(\words[14]/data_i[13] ) );
  AO22X1 U4426 ( .IN1(\read_value_mux[14][14] ), .IN2(n1624), .IN3(
        write_data[14]), .IN4(n3147), .Q(\words[14]/data_i[14] ) );
  AO22X1 U4427 ( .IN1(\read_value_mux[14][15] ), .IN2(n1624), .IN3(
        write_data[15]), .IN4(n3147), .Q(\words[14]/data_i[15] ) );
  AO22X1 U4428 ( .IN1(\read_value_mux[14][16] ), .IN2(n1624), .IN3(
        write_data[16]), .IN4(n3147), .Q(\words[14]/data_i[16] ) );
  AO22X1 U4429 ( .IN1(\read_value_mux[14][17] ), .IN2(n1624), .IN3(
        write_data[17]), .IN4(n3147), .Q(\words[14]/data_i[17] ) );
  AO22X1 U4430 ( .IN1(\read_value_mux[14][18] ), .IN2(n1624), .IN3(
        write_data[18]), .IN4(n3147), .Q(\words[14]/data_i[18] ) );
  AO22X1 U4431 ( .IN1(\read_value_mux[14][19] ), .IN2(n1624), .IN3(
        write_data[19]), .IN4(n3147), .Q(\words[14]/data_i[19] ) );
  AO22X1 U4432 ( .IN1(\read_value_mux[14][1] ), .IN2(n1624), .IN3(
        write_data[1]), .IN4(n3147), .Q(\words[14]/data_i[1] ) );
  AO22X1 U4433 ( .IN1(\read_value_mux[14][20] ), .IN2(n1624), .IN3(
        write_data[20]), .IN4(n3147), .Q(\words[14]/data_i[20] ) );
  AO22X1 U4434 ( .IN1(\read_value_mux[14][21] ), .IN2(n1624), .IN3(
        write_data[21]), .IN4(n3147), .Q(\words[14]/data_i[21] ) );
  AO22X1 U4435 ( .IN1(\read_value_mux[14][22] ), .IN2(n1624), .IN3(
        write_data[22]), .IN4(n3147), .Q(\words[14]/data_i[22] ) );
  AO22X1 U4436 ( .IN1(\read_value_mux[14][23] ), .IN2(n1624), .IN3(
        write_data[23]), .IN4(n3147), .Q(\words[14]/data_i[23] ) );
  AO22X1 U4437 ( .IN1(\read_value_mux[14][24] ), .IN2(n1624), .IN3(
        write_data[24]), .IN4(n3147), .Q(\words[14]/data_i[24] ) );
  AO22X1 U4438 ( .IN1(\read_value_mux[14][25] ), .IN2(n1624), .IN3(
        write_data[25]), .IN4(n3147), .Q(\words[14]/data_i[25] ) );
  AO22X1 U4439 ( .IN1(\read_value_mux[14][26] ), .IN2(n1624), .IN3(
        write_data[26]), .IN4(n3147), .Q(\words[14]/data_i[26] ) );
  AO22X1 U4440 ( .IN1(\read_value_mux[14][27] ), .IN2(n1624), .IN3(
        write_data[27]), .IN4(n3147), .Q(\words[14]/data_i[27] ) );
  AO22X1 U4441 ( .IN1(\read_value_mux[14][28] ), .IN2(n1624), .IN3(
        write_data[28]), .IN4(n3147), .Q(\words[14]/data_i[28] ) );
  AO22X1 U4442 ( .IN1(\read_value_mux[14][29] ), .IN2(n1624), .IN3(
        write_data[29]), .IN4(n3147), .Q(\words[14]/data_i[29] ) );
  AO22X1 U4443 ( .IN1(\read_value_mux[14][2] ), .IN2(n1624), .IN3(
        write_data[2]), .IN4(n3147), .Q(\words[14]/data_i[2] ) );
  AO22X1 U4444 ( .IN1(\read_value_mux[14][30] ), .IN2(n1624), .IN3(
        write_data[30]), .IN4(n3147), .Q(\words[14]/data_i[30] ) );
  AO22X1 U4445 ( .IN1(\read_value_mux[14][31] ), .IN2(n1624), .IN3(
        write_data[31]), .IN4(n3147), .Q(\words[14]/data_i[31] ) );
  AO22X1 U4446 ( .IN1(\read_value_mux[14][3] ), .IN2(n1624), .IN3(
        write_data[3]), .IN4(n3147), .Q(\words[14]/data_i[3] ) );
  AO22X1 U4447 ( .IN1(\read_value_mux[14][4] ), .IN2(n1624), .IN3(
        write_data[4]), .IN4(n3147), .Q(\words[14]/data_i[4] ) );
  AO22X1 U4448 ( .IN1(\read_value_mux[14][5] ), .IN2(n1624), .IN3(
        write_data[5]), .IN4(n3147), .Q(\words[14]/data_i[5] ) );
  AO22X1 U4449 ( .IN1(\read_value_mux[14][6] ), .IN2(n1624), .IN3(
        write_data[6]), .IN4(n3147), .Q(\words[14]/data_i[6] ) );
  AO22X1 U4450 ( .IN1(\read_value_mux[14][7] ), .IN2(n1624), .IN3(
        write_data[7]), .IN4(n3147), .Q(\words[14]/data_i[7] ) );
  AO22X1 U4451 ( .IN1(\read_value_mux[14][8] ), .IN2(n1624), .IN3(
        write_data[8]), .IN4(n3147), .Q(\words[14]/data_i[8] ) );
  AO22X1 U4452 ( .IN1(\read_value_mux[14][9] ), .IN2(n1624), .IN3(
        write_data[9]), .IN4(n3147), .Q(\words[14]/data_i[9] ) );
  AO21X1 U4453 ( .IN1(\words[14]/valid_o ), .IN2(n1743), .IN3(n3147), .Q(
        \words[14]/valid_i ) );
  AO22X1 U4454 ( .IN1(\read_value_mux[15][0] ), .IN2(n1625), .IN3(
        write_data[0]), .IN4(n3149), .Q(\words[15]/data_i[0] ) );
  AO22X1 U4455 ( .IN1(\read_value_mux[15][10] ), .IN2(n1625), .IN3(
        write_data[10]), .IN4(n3149), .Q(\words[15]/data_i[10] ) );
  AO22X1 U4456 ( .IN1(\read_value_mux[15][11] ), .IN2(n1625), .IN3(
        write_data[11]), .IN4(n3149), .Q(\words[15]/data_i[11] ) );
  AO22X1 U4457 ( .IN1(\read_value_mux[15][12] ), .IN2(n1625), .IN3(
        write_data[12]), .IN4(n3149), .Q(\words[15]/data_i[12] ) );
  AO22X1 U4458 ( .IN1(\read_value_mux[15][13] ), .IN2(n1625), .IN3(
        write_data[13]), .IN4(n3149), .Q(\words[15]/data_i[13] ) );
  AO22X1 U4459 ( .IN1(\read_value_mux[15][14] ), .IN2(n1625), .IN3(
        write_data[14]), .IN4(n3149), .Q(\words[15]/data_i[14] ) );
  AO22X1 U4460 ( .IN1(\read_value_mux[15][15] ), .IN2(n1625), .IN3(
        write_data[15]), .IN4(n3149), .Q(\words[15]/data_i[15] ) );
  AO22X1 U4461 ( .IN1(\read_value_mux[15][16] ), .IN2(n1625), .IN3(
        write_data[16]), .IN4(n3149), .Q(\words[15]/data_i[16] ) );
  AO22X1 U4462 ( .IN1(\read_value_mux[15][17] ), .IN2(n1625), .IN3(
        write_data[17]), .IN4(n3149), .Q(\words[15]/data_i[17] ) );
  AO22X1 U4463 ( .IN1(\read_value_mux[15][18] ), .IN2(n1625), .IN3(
        write_data[18]), .IN4(n3149), .Q(\words[15]/data_i[18] ) );
  AO22X1 U4464 ( .IN1(\read_value_mux[15][19] ), .IN2(n1625), .IN3(
        write_data[19]), .IN4(n3149), .Q(\words[15]/data_i[19] ) );
  AO22X1 U4465 ( .IN1(\read_value_mux[15][1] ), .IN2(n1625), .IN3(
        write_data[1]), .IN4(n3149), .Q(\words[15]/data_i[1] ) );
  AO22X1 U4466 ( .IN1(\read_value_mux[15][20] ), .IN2(n1625), .IN3(
        write_data[20]), .IN4(n3149), .Q(\words[15]/data_i[20] ) );
  AO22X1 U4467 ( .IN1(\read_value_mux[15][21] ), .IN2(n1625), .IN3(
        write_data[21]), .IN4(n3149), .Q(\words[15]/data_i[21] ) );
  AO22X1 U4468 ( .IN1(\read_value_mux[15][22] ), .IN2(n1625), .IN3(
        write_data[22]), .IN4(n3149), .Q(\words[15]/data_i[22] ) );
  AO22X1 U4469 ( .IN1(\read_value_mux[15][23] ), .IN2(n1625), .IN3(
        write_data[23]), .IN4(n3149), .Q(\words[15]/data_i[23] ) );
  AO22X1 U4470 ( .IN1(\read_value_mux[15][24] ), .IN2(n1625), .IN3(
        write_data[24]), .IN4(n3149), .Q(\words[15]/data_i[24] ) );
  AO22X1 U4471 ( .IN1(\read_value_mux[15][25] ), .IN2(n1625), .IN3(
        write_data[25]), .IN4(n3149), .Q(\words[15]/data_i[25] ) );
  AO22X1 U4472 ( .IN1(\read_value_mux[15][26] ), .IN2(n1625), .IN3(
        write_data[26]), .IN4(n3149), .Q(\words[15]/data_i[26] ) );
  AO22X1 U4473 ( .IN1(\read_value_mux[15][27] ), .IN2(n1625), .IN3(
        write_data[27]), .IN4(n3149), .Q(\words[15]/data_i[27] ) );
  AO22X1 U4474 ( .IN1(\read_value_mux[15][28] ), .IN2(n1625), .IN3(
        write_data[28]), .IN4(n3149), .Q(\words[15]/data_i[28] ) );
  AO22X1 U4475 ( .IN1(\read_value_mux[15][29] ), .IN2(n1625), .IN3(
        write_data[29]), .IN4(n3149), .Q(\words[15]/data_i[29] ) );
  AO22X1 U4476 ( .IN1(\read_value_mux[15][2] ), .IN2(n1625), .IN3(
        write_data[2]), .IN4(n3149), .Q(\words[15]/data_i[2] ) );
  AO22X1 U4477 ( .IN1(\read_value_mux[15][30] ), .IN2(n1625), .IN3(
        write_data[30]), .IN4(n3149), .Q(\words[15]/data_i[30] ) );
  AO22X1 U4478 ( .IN1(\read_value_mux[15][31] ), .IN2(n1625), .IN3(
        write_data[31]), .IN4(n3149), .Q(\words[15]/data_i[31] ) );
  AO22X1 U4479 ( .IN1(\read_value_mux[15][3] ), .IN2(n1625), .IN3(
        write_data[3]), .IN4(n3149), .Q(\words[15]/data_i[3] ) );
  AO22X1 U4480 ( .IN1(\read_value_mux[15][4] ), .IN2(n1625), .IN3(
        write_data[4]), .IN4(n3149), .Q(\words[15]/data_i[4] ) );
  AO22X1 U4481 ( .IN1(\read_value_mux[15][5] ), .IN2(n1625), .IN3(
        write_data[5]), .IN4(n3149), .Q(\words[15]/data_i[5] ) );
  AO22X1 U4482 ( .IN1(\read_value_mux[15][6] ), .IN2(n1625), .IN3(
        write_data[6]), .IN4(n3149), .Q(\words[15]/data_i[6] ) );
  AO22X1 U4483 ( .IN1(\read_value_mux[15][7] ), .IN2(n1625), .IN3(
        write_data[7]), .IN4(n3149), .Q(\words[15]/data_i[7] ) );
  AO22X1 U4484 ( .IN1(\read_value_mux[15][8] ), .IN2(n1625), .IN3(
        write_data[8]), .IN4(n3149), .Q(\words[15]/data_i[8] ) );
  AO22X1 U4485 ( .IN1(\read_value_mux[15][9] ), .IN2(n1625), .IN3(
        write_data[9]), .IN4(n3149), .Q(\words[15]/data_i[9] ) );
  AO21X1 U4486 ( .IN1(\words[15]/valid_o ), .IN2(n1743), .IN3(n3149), .Q(
        \words[15]/valid_i ) );
  AO22X1 U4487 ( .IN1(\read_value_mux[16][0] ), .IN2(n1620), .IN3(
        write_data[0]), .IN4(n3153), .Q(\words[16]/data_i[0] ) );
  AO22X1 U4488 ( .IN1(\read_value_mux[16][10] ), .IN2(n1620), .IN3(
        write_data[10]), .IN4(n3153), .Q(\words[16]/data_i[10] ) );
  AO22X1 U4489 ( .IN1(\read_value_mux[16][11] ), .IN2(n1620), .IN3(
        write_data[11]), .IN4(n3153), .Q(\words[16]/data_i[11] ) );
  AO22X1 U4490 ( .IN1(\read_value_mux[16][12] ), .IN2(n1620), .IN3(
        write_data[12]), .IN4(n3153), .Q(\words[16]/data_i[12] ) );
  AO22X1 U4491 ( .IN1(\read_value_mux[16][13] ), .IN2(n1620), .IN3(
        write_data[13]), .IN4(n3153), .Q(\words[16]/data_i[13] ) );
  AO22X1 U4492 ( .IN1(\read_value_mux[16][14] ), .IN2(n1620), .IN3(
        write_data[14]), .IN4(n3153), .Q(\words[16]/data_i[14] ) );
  AO22X1 U4493 ( .IN1(\read_value_mux[16][15] ), .IN2(n1620), .IN3(
        write_data[15]), .IN4(n3153), .Q(\words[16]/data_i[15] ) );
  AO22X1 U4494 ( .IN1(\read_value_mux[16][16] ), .IN2(n1620), .IN3(
        write_data[16]), .IN4(n3153), .Q(\words[16]/data_i[16] ) );
  AO22X1 U4495 ( .IN1(\read_value_mux[16][17] ), .IN2(n1620), .IN3(
        write_data[17]), .IN4(n3153), .Q(\words[16]/data_i[17] ) );
  AO22X1 U4496 ( .IN1(\read_value_mux[16][18] ), .IN2(n1620), .IN3(
        write_data[18]), .IN4(n3153), .Q(\words[16]/data_i[18] ) );
  AO22X1 U4497 ( .IN1(\read_value_mux[16][19] ), .IN2(n1620), .IN3(
        write_data[19]), .IN4(n3153), .Q(\words[16]/data_i[19] ) );
  AO22X1 U4498 ( .IN1(\read_value_mux[16][1] ), .IN2(n1620), .IN3(
        write_data[1]), .IN4(n3153), .Q(\words[16]/data_i[1] ) );
  AO22X1 U4499 ( .IN1(\read_value_mux[16][20] ), .IN2(n1620), .IN3(
        write_data[20]), .IN4(n3153), .Q(\words[16]/data_i[20] ) );
  AO22X1 U4500 ( .IN1(\read_value_mux[16][21] ), .IN2(n1620), .IN3(
        write_data[21]), .IN4(n3153), .Q(\words[16]/data_i[21] ) );
  AO22X1 U4501 ( .IN1(\read_value_mux[16][22] ), .IN2(n1620), .IN3(
        write_data[22]), .IN4(n3153), .Q(\words[16]/data_i[22] ) );
  AO22X1 U4502 ( .IN1(\read_value_mux[16][23] ), .IN2(n1620), .IN3(
        write_data[23]), .IN4(n3153), .Q(\words[16]/data_i[23] ) );
  AO22X1 U4503 ( .IN1(\read_value_mux[16][24] ), .IN2(n1620), .IN3(
        write_data[24]), .IN4(n3153), .Q(\words[16]/data_i[24] ) );
  AO22X1 U4504 ( .IN1(\read_value_mux[16][25] ), .IN2(n1620), .IN3(
        write_data[25]), .IN4(n3153), .Q(\words[16]/data_i[25] ) );
  AO22X1 U4505 ( .IN1(\read_value_mux[16][26] ), .IN2(n1620), .IN3(
        write_data[26]), .IN4(n3153), .Q(\words[16]/data_i[26] ) );
  AO22X1 U4506 ( .IN1(\read_value_mux[16][27] ), .IN2(n1620), .IN3(
        write_data[27]), .IN4(n3153), .Q(\words[16]/data_i[27] ) );
  AO22X1 U4507 ( .IN1(\read_value_mux[16][28] ), .IN2(n1620), .IN3(
        write_data[28]), .IN4(n3153), .Q(\words[16]/data_i[28] ) );
  AO22X1 U4508 ( .IN1(\read_value_mux[16][29] ), .IN2(n1620), .IN3(
        write_data[29]), .IN4(n3153), .Q(\words[16]/data_i[29] ) );
  AO22X1 U4509 ( .IN1(\read_value_mux[16][2] ), .IN2(n1620), .IN3(
        write_data[2]), .IN4(n3153), .Q(\words[16]/data_i[2] ) );
  AO22X1 U4510 ( .IN1(\read_value_mux[16][30] ), .IN2(n1620), .IN3(
        write_data[30]), .IN4(n3153), .Q(\words[16]/data_i[30] ) );
  AO22X1 U4511 ( .IN1(\read_value_mux[16][31] ), .IN2(n1620), .IN3(
        write_data[31]), .IN4(n3153), .Q(\words[16]/data_i[31] ) );
  AO22X1 U4512 ( .IN1(\read_value_mux[16][3] ), .IN2(n1620), .IN3(
        write_data[3]), .IN4(n3153), .Q(\words[16]/data_i[3] ) );
  AO22X1 U4513 ( .IN1(\read_value_mux[16][4] ), .IN2(n1620), .IN3(
        write_data[4]), .IN4(n3153), .Q(\words[16]/data_i[4] ) );
  AO22X1 U4514 ( .IN1(\read_value_mux[16][5] ), .IN2(n1620), .IN3(
        write_data[5]), .IN4(n3153), .Q(\words[16]/data_i[5] ) );
  AO22X1 U4515 ( .IN1(\read_value_mux[16][6] ), .IN2(n1620), .IN3(
        write_data[6]), .IN4(n3153), .Q(\words[16]/data_i[6] ) );
  AO22X1 U4516 ( .IN1(\read_value_mux[16][7] ), .IN2(n1620), .IN3(
        write_data[7]), .IN4(n3153), .Q(\words[16]/data_i[7] ) );
  AO22X1 U4517 ( .IN1(\read_value_mux[16][8] ), .IN2(n1620), .IN3(
        write_data[8]), .IN4(n3153), .Q(\words[16]/data_i[8] ) );
  AO22X1 U4518 ( .IN1(\read_value_mux[16][9] ), .IN2(n1620), .IN3(
        write_data[9]), .IN4(n3153), .Q(\words[16]/data_i[9] ) );
  AO21X1 U4519 ( .IN1(\words[16]/valid_o ), .IN2(n1743), .IN3(n3153), .Q(
        \words[16]/valid_i ) );
  AO22X1 U4520 ( .IN1(\read_value_mux[17][0] ), .IN2(n1621), .IN3(
        write_data[0]), .IN4(n3154), .Q(\words[17]/data_i[0] ) );
  AO22X1 U4521 ( .IN1(\read_value_mux[17][10] ), .IN2(n1621), .IN3(
        write_data[10]), .IN4(n3154), .Q(\words[17]/data_i[10] ) );
  AO22X1 U4522 ( .IN1(\read_value_mux[17][11] ), .IN2(n1621), .IN3(
        write_data[11]), .IN4(n3154), .Q(\words[17]/data_i[11] ) );
  AO22X1 U4523 ( .IN1(\read_value_mux[17][12] ), .IN2(n1621), .IN3(
        write_data[12]), .IN4(n3154), .Q(\words[17]/data_i[12] ) );
  AO22X1 U4524 ( .IN1(\read_value_mux[17][13] ), .IN2(n1621), .IN3(
        write_data[13]), .IN4(n3154), .Q(\words[17]/data_i[13] ) );
  AO22X1 U4525 ( .IN1(\read_value_mux[17][14] ), .IN2(n1621), .IN3(
        write_data[14]), .IN4(n3154), .Q(\words[17]/data_i[14] ) );
  AO22X1 U4526 ( .IN1(\read_value_mux[17][15] ), .IN2(n1621), .IN3(
        write_data[15]), .IN4(n3154), .Q(\words[17]/data_i[15] ) );
  AO22X1 U4527 ( .IN1(\read_value_mux[17][16] ), .IN2(n1621), .IN3(
        write_data[16]), .IN4(n3154), .Q(\words[17]/data_i[16] ) );
  AO22X1 U4528 ( .IN1(\read_value_mux[17][17] ), .IN2(n1621), .IN3(
        write_data[17]), .IN4(n3154), .Q(\words[17]/data_i[17] ) );
  AO22X1 U4529 ( .IN1(\read_value_mux[17][18] ), .IN2(n1621), .IN3(
        write_data[18]), .IN4(n3154), .Q(\words[17]/data_i[18] ) );
  AO22X1 U4530 ( .IN1(\read_value_mux[17][19] ), .IN2(n1621), .IN3(
        write_data[19]), .IN4(n3154), .Q(\words[17]/data_i[19] ) );
  AO22X1 U4531 ( .IN1(\read_value_mux[17][1] ), .IN2(n1621), .IN3(
        write_data[1]), .IN4(n3154), .Q(\words[17]/data_i[1] ) );
  AO22X1 U4532 ( .IN1(\read_value_mux[17][20] ), .IN2(n1621), .IN3(
        write_data[20]), .IN4(n3154), .Q(\words[17]/data_i[20] ) );
  AO22X1 U4533 ( .IN1(\read_value_mux[17][21] ), .IN2(n1621), .IN3(
        write_data[21]), .IN4(n3154), .Q(\words[17]/data_i[21] ) );
  AO22X1 U4534 ( .IN1(\read_value_mux[17][22] ), .IN2(n1621), .IN3(
        write_data[22]), .IN4(n3154), .Q(\words[17]/data_i[22] ) );
  AO22X1 U4535 ( .IN1(\read_value_mux[17][23] ), .IN2(n1621), .IN3(
        write_data[23]), .IN4(n3154), .Q(\words[17]/data_i[23] ) );
  AO22X1 U4536 ( .IN1(\read_value_mux[17][24] ), .IN2(n1621), .IN3(
        write_data[24]), .IN4(n3154), .Q(\words[17]/data_i[24] ) );
  AO22X1 U4537 ( .IN1(\read_value_mux[17][25] ), .IN2(n1621), .IN3(
        write_data[25]), .IN4(n3154), .Q(\words[17]/data_i[25] ) );
  AO22X1 U4538 ( .IN1(\read_value_mux[17][26] ), .IN2(n1621), .IN3(
        write_data[26]), .IN4(n3154), .Q(\words[17]/data_i[26] ) );
  AO22X1 U4539 ( .IN1(\read_value_mux[17][27] ), .IN2(n1621), .IN3(
        write_data[27]), .IN4(n3154), .Q(\words[17]/data_i[27] ) );
  AO22X1 U4540 ( .IN1(\read_value_mux[17][28] ), .IN2(n1621), .IN3(
        write_data[28]), .IN4(n3154), .Q(\words[17]/data_i[28] ) );
  AO22X1 U4541 ( .IN1(\read_value_mux[17][29] ), .IN2(n1621), .IN3(
        write_data[29]), .IN4(n3154), .Q(\words[17]/data_i[29] ) );
  AO22X1 U4542 ( .IN1(\read_value_mux[17][2] ), .IN2(n1621), .IN3(
        write_data[2]), .IN4(n3154), .Q(\words[17]/data_i[2] ) );
  AO22X1 U4543 ( .IN1(\read_value_mux[17][30] ), .IN2(n1621), .IN3(
        write_data[30]), .IN4(n3154), .Q(\words[17]/data_i[30] ) );
  AO22X1 U4544 ( .IN1(\read_value_mux[17][31] ), .IN2(n1621), .IN3(
        write_data[31]), .IN4(n3154), .Q(\words[17]/data_i[31] ) );
  AO22X1 U4545 ( .IN1(\read_value_mux[17][3] ), .IN2(n1621), .IN3(
        write_data[3]), .IN4(n3154), .Q(\words[17]/data_i[3] ) );
  AO22X1 U4546 ( .IN1(\read_value_mux[17][4] ), .IN2(n1621), .IN3(
        write_data[4]), .IN4(n3154), .Q(\words[17]/data_i[4] ) );
  AO22X1 U4547 ( .IN1(\read_value_mux[17][5] ), .IN2(n1621), .IN3(
        write_data[5]), .IN4(n3154), .Q(\words[17]/data_i[5] ) );
  AO22X1 U4548 ( .IN1(\read_value_mux[17][6] ), .IN2(n1621), .IN3(
        write_data[6]), .IN4(n3154), .Q(\words[17]/data_i[6] ) );
  AO22X1 U4549 ( .IN1(\read_value_mux[17][7] ), .IN2(n1621), .IN3(
        write_data[7]), .IN4(n3154), .Q(\words[17]/data_i[7] ) );
  AO22X1 U4550 ( .IN1(\read_value_mux[17][8] ), .IN2(n1621), .IN3(
        write_data[8]), .IN4(n3154), .Q(\words[17]/data_i[8] ) );
  AO22X1 U4551 ( .IN1(\read_value_mux[17][9] ), .IN2(n1621), .IN3(
        write_data[9]), .IN4(n3154), .Q(\words[17]/data_i[9] ) );
  AO21X1 U4552 ( .IN1(\words[17]/valid_o ), .IN2(n1743), .IN3(n3154), .Q(
        \words[17]/valid_i ) );
  AO22X1 U4553 ( .IN1(\read_value_mux[18][0] ), .IN2(n1626), .IN3(
        write_data[0]), .IN4(n3155), .Q(\words[18]/data_i[0] ) );
  AO22X1 U4554 ( .IN1(\read_value_mux[18][10] ), .IN2(n1626), .IN3(
        write_data[10]), .IN4(n3155), .Q(\words[18]/data_i[10] ) );
  AO22X1 U4555 ( .IN1(\read_value_mux[18][11] ), .IN2(n1626), .IN3(
        write_data[11]), .IN4(n3155), .Q(\words[18]/data_i[11] ) );
  AO22X1 U4556 ( .IN1(\read_value_mux[18][12] ), .IN2(n1626), .IN3(
        write_data[12]), .IN4(n3155), .Q(\words[18]/data_i[12] ) );
  AO22X1 U4557 ( .IN1(\read_value_mux[18][13] ), .IN2(n1626), .IN3(
        write_data[13]), .IN4(n3155), .Q(\words[18]/data_i[13] ) );
  AO22X1 U4558 ( .IN1(\read_value_mux[18][14] ), .IN2(n1626), .IN3(
        write_data[14]), .IN4(n3155), .Q(\words[18]/data_i[14] ) );
  AO22X1 U4559 ( .IN1(\read_value_mux[18][15] ), .IN2(n1626), .IN3(
        write_data[15]), .IN4(n3155), .Q(\words[18]/data_i[15] ) );
  AO22X1 U4560 ( .IN1(\read_value_mux[18][16] ), .IN2(n1626), .IN3(
        write_data[16]), .IN4(n3155), .Q(\words[18]/data_i[16] ) );
  AO22X1 U4561 ( .IN1(\read_value_mux[18][17] ), .IN2(n1626), .IN3(
        write_data[17]), .IN4(n3155), .Q(\words[18]/data_i[17] ) );
  AO22X1 U4562 ( .IN1(\read_value_mux[18][18] ), .IN2(n1626), .IN3(
        write_data[18]), .IN4(n3155), .Q(\words[18]/data_i[18] ) );
  AO22X1 U4563 ( .IN1(\read_value_mux[18][19] ), .IN2(n1626), .IN3(
        write_data[19]), .IN4(n3155), .Q(\words[18]/data_i[19] ) );
  AO22X1 U4564 ( .IN1(\read_value_mux[18][1] ), .IN2(n1626), .IN3(
        write_data[1]), .IN4(n3155), .Q(\words[18]/data_i[1] ) );
  AO22X1 U4565 ( .IN1(\read_value_mux[18][20] ), .IN2(n1626), .IN3(
        write_data[20]), .IN4(n3155), .Q(\words[18]/data_i[20] ) );
  AO22X1 U4566 ( .IN1(\read_value_mux[18][21] ), .IN2(n1626), .IN3(
        write_data[21]), .IN4(n3155), .Q(\words[18]/data_i[21] ) );
  AO22X1 U4567 ( .IN1(\read_value_mux[18][22] ), .IN2(n1626), .IN3(
        write_data[22]), .IN4(n3155), .Q(\words[18]/data_i[22] ) );
  AO22X1 U4568 ( .IN1(\read_value_mux[18][23] ), .IN2(n1626), .IN3(
        write_data[23]), .IN4(n3155), .Q(\words[18]/data_i[23] ) );
  AO22X1 U4569 ( .IN1(\read_value_mux[18][24] ), .IN2(n1626), .IN3(
        write_data[24]), .IN4(n3155), .Q(\words[18]/data_i[24] ) );
  AO22X1 U4570 ( .IN1(\read_value_mux[18][25] ), .IN2(n1626), .IN3(
        write_data[25]), .IN4(n3155), .Q(\words[18]/data_i[25] ) );
  AO22X1 U4571 ( .IN1(\read_value_mux[18][26] ), .IN2(n1626), .IN3(
        write_data[26]), .IN4(n3155), .Q(\words[18]/data_i[26] ) );
  AO22X1 U4572 ( .IN1(\read_value_mux[18][27] ), .IN2(n1626), .IN3(
        write_data[27]), .IN4(n3155), .Q(\words[18]/data_i[27] ) );
  AO22X1 U4573 ( .IN1(\read_value_mux[18][28] ), .IN2(n1626), .IN3(
        write_data[28]), .IN4(n3155), .Q(\words[18]/data_i[28] ) );
  AO22X1 U4574 ( .IN1(\read_value_mux[18][29] ), .IN2(n1626), .IN3(
        write_data[29]), .IN4(n3155), .Q(\words[18]/data_i[29] ) );
  AO22X1 U4575 ( .IN1(\read_value_mux[18][2] ), .IN2(n1626), .IN3(
        write_data[2]), .IN4(n3155), .Q(\words[18]/data_i[2] ) );
  AO22X1 U4576 ( .IN1(\read_value_mux[18][30] ), .IN2(n1626), .IN3(
        write_data[30]), .IN4(n3155), .Q(\words[18]/data_i[30] ) );
  AO22X1 U4577 ( .IN1(\read_value_mux[18][31] ), .IN2(n1626), .IN3(
        write_data[31]), .IN4(n3155), .Q(\words[18]/data_i[31] ) );
  AO22X1 U4578 ( .IN1(\read_value_mux[18][3] ), .IN2(n1626), .IN3(
        write_data[3]), .IN4(n3155), .Q(\words[18]/data_i[3] ) );
  AO22X1 U4579 ( .IN1(\read_value_mux[18][4] ), .IN2(n1626), .IN3(
        write_data[4]), .IN4(n3155), .Q(\words[18]/data_i[4] ) );
  AO22X1 U4580 ( .IN1(\read_value_mux[18][5] ), .IN2(n1626), .IN3(
        write_data[5]), .IN4(n3155), .Q(\words[18]/data_i[5] ) );
  AO22X1 U4581 ( .IN1(\read_value_mux[18][6] ), .IN2(n1626), .IN3(
        write_data[6]), .IN4(n3155), .Q(\words[18]/data_i[6] ) );
  AO22X1 U4582 ( .IN1(\read_value_mux[18][7] ), .IN2(n1626), .IN3(
        write_data[7]), .IN4(n3155), .Q(\words[18]/data_i[7] ) );
  AO22X1 U4583 ( .IN1(\read_value_mux[18][8] ), .IN2(n1626), .IN3(
        write_data[8]), .IN4(n3155), .Q(\words[18]/data_i[8] ) );
  AO22X1 U4584 ( .IN1(\read_value_mux[18][9] ), .IN2(n1626), .IN3(
        write_data[9]), .IN4(n3155), .Q(\words[18]/data_i[9] ) );
  AO21X1 U4585 ( .IN1(\words[18]/valid_o ), .IN2(n1743), .IN3(n3155), .Q(
        \words[18]/valid_i ) );
  AO22X1 U4586 ( .IN1(\read_value_mux[19][0] ), .IN2(n1627), .IN3(
        write_data[0]), .IN4(n3157), .Q(\words[19]/data_i[0] ) );
  AO22X1 U4587 ( .IN1(\read_value_mux[19][10] ), .IN2(n1627), .IN3(
        write_data[10]), .IN4(n3157), .Q(\words[19]/data_i[10] ) );
  AO22X1 U4588 ( .IN1(\read_value_mux[19][11] ), .IN2(n1627), .IN3(
        write_data[11]), .IN4(n3157), .Q(\words[19]/data_i[11] ) );
  AO22X1 U4589 ( .IN1(\read_value_mux[19][12] ), .IN2(n1627), .IN3(
        write_data[12]), .IN4(n3157), .Q(\words[19]/data_i[12] ) );
  AO22X1 U4590 ( .IN1(\read_value_mux[19][13] ), .IN2(n1627), .IN3(
        write_data[13]), .IN4(n3157), .Q(\words[19]/data_i[13] ) );
  AO22X1 U4591 ( .IN1(\read_value_mux[19][14] ), .IN2(n1627), .IN3(
        write_data[14]), .IN4(n3157), .Q(\words[19]/data_i[14] ) );
  AO22X1 U4592 ( .IN1(\read_value_mux[19][15] ), .IN2(n1627), .IN3(
        write_data[15]), .IN4(n3157), .Q(\words[19]/data_i[15] ) );
  AO22X1 U4593 ( .IN1(\read_value_mux[19][16] ), .IN2(n1627), .IN3(
        write_data[16]), .IN4(n3157), .Q(\words[19]/data_i[16] ) );
  AO22X1 U4594 ( .IN1(\read_value_mux[19][17] ), .IN2(n1627), .IN3(
        write_data[17]), .IN4(n3157), .Q(\words[19]/data_i[17] ) );
  AO22X1 U4595 ( .IN1(\read_value_mux[19][18] ), .IN2(n1627), .IN3(
        write_data[18]), .IN4(n3157), .Q(\words[19]/data_i[18] ) );
  AO22X1 U4596 ( .IN1(\read_value_mux[19][19] ), .IN2(n1627), .IN3(
        write_data[19]), .IN4(n3157), .Q(\words[19]/data_i[19] ) );
  AO22X1 U4597 ( .IN1(\read_value_mux[19][1] ), .IN2(n1627), .IN3(
        write_data[1]), .IN4(n3157), .Q(\words[19]/data_i[1] ) );
  AO22X1 U4598 ( .IN1(\read_value_mux[19][20] ), .IN2(n1627), .IN3(
        write_data[20]), .IN4(n3157), .Q(\words[19]/data_i[20] ) );
  AO22X1 U4599 ( .IN1(\read_value_mux[19][21] ), .IN2(n1627), .IN3(
        write_data[21]), .IN4(n3157), .Q(\words[19]/data_i[21] ) );
  AO22X1 U4600 ( .IN1(\read_value_mux[19][22] ), .IN2(n1627), .IN3(
        write_data[22]), .IN4(n3157), .Q(\words[19]/data_i[22] ) );
  AO22X1 U4601 ( .IN1(\read_value_mux[19][23] ), .IN2(n1627), .IN3(
        write_data[23]), .IN4(n3157), .Q(\words[19]/data_i[23] ) );
  AO22X1 U4602 ( .IN1(\read_value_mux[19][24] ), .IN2(n1627), .IN3(
        write_data[24]), .IN4(n3157), .Q(\words[19]/data_i[24] ) );
  AO22X1 U4603 ( .IN1(\read_value_mux[19][25] ), .IN2(n1627), .IN3(
        write_data[25]), .IN4(n3157), .Q(\words[19]/data_i[25] ) );
  AO22X1 U4604 ( .IN1(\read_value_mux[19][26] ), .IN2(n1627), .IN3(
        write_data[26]), .IN4(n3157), .Q(\words[19]/data_i[26] ) );
  AO22X1 U4605 ( .IN1(\read_value_mux[19][27] ), .IN2(n1627), .IN3(
        write_data[27]), .IN4(n3157), .Q(\words[19]/data_i[27] ) );
  AO22X1 U4606 ( .IN1(\read_value_mux[19][28] ), .IN2(n1627), .IN3(
        write_data[28]), .IN4(n3157), .Q(\words[19]/data_i[28] ) );
  AO22X1 U4607 ( .IN1(\read_value_mux[19][29] ), .IN2(n1627), .IN3(
        write_data[29]), .IN4(n3157), .Q(\words[19]/data_i[29] ) );
  AO22X1 U4608 ( .IN1(\read_value_mux[19][2] ), .IN2(n1627), .IN3(
        write_data[2]), .IN4(n3157), .Q(\words[19]/data_i[2] ) );
  AO22X1 U4609 ( .IN1(\read_value_mux[19][30] ), .IN2(n1627), .IN3(
        write_data[30]), .IN4(n3157), .Q(\words[19]/data_i[30] ) );
  AO22X1 U4610 ( .IN1(\read_value_mux[19][31] ), .IN2(n1627), .IN3(
        write_data[31]), .IN4(n3157), .Q(\words[19]/data_i[31] ) );
  AO22X1 U4611 ( .IN1(\read_value_mux[19][3] ), .IN2(n1627), .IN3(
        write_data[3]), .IN4(n3157), .Q(\words[19]/data_i[3] ) );
  AO22X1 U4612 ( .IN1(\read_value_mux[19][4] ), .IN2(n1627), .IN3(
        write_data[4]), .IN4(n3157), .Q(\words[19]/data_i[4] ) );
  AO22X1 U4613 ( .IN1(\read_value_mux[19][5] ), .IN2(n1627), .IN3(
        write_data[5]), .IN4(n3157), .Q(\words[19]/data_i[5] ) );
  AO22X1 U4614 ( .IN1(\read_value_mux[19][6] ), .IN2(n1627), .IN3(
        write_data[6]), .IN4(n3157), .Q(\words[19]/data_i[6] ) );
  AO22X1 U4615 ( .IN1(\read_value_mux[19][7] ), .IN2(n1627), .IN3(
        write_data[7]), .IN4(n3157), .Q(\words[19]/data_i[7] ) );
  AO22X1 U4616 ( .IN1(\read_value_mux[19][8] ), .IN2(n1627), .IN3(
        write_data[8]), .IN4(n3157), .Q(\words[19]/data_i[8] ) );
  AO22X1 U4617 ( .IN1(\read_value_mux[19][9] ), .IN2(n1627), .IN3(
        write_data[9]), .IN4(n3157), .Q(\words[19]/data_i[9] ) );
  AO21X1 U4618 ( .IN1(\words[19]/valid_o ), .IN2(n1743), .IN3(n3157), .Q(
        \words[19]/valid_i ) );
  AO22X1 U4619 ( .IN1(\read_value_mux[1][0] ), .IN2(n1622), .IN3(write_data[0]), .IN4(n3158), .Q(\words[1]/data_i[0] ) );
  AO22X1 U4620 ( .IN1(\read_value_mux[1][10] ), .IN2(n1622), .IN3(
        write_data[10]), .IN4(n3158), .Q(\words[1]/data_i[10] ) );
  AO22X1 U4621 ( .IN1(\read_value_mux[1][11] ), .IN2(n1622), .IN3(
        write_data[11]), .IN4(n3158), .Q(\words[1]/data_i[11] ) );
  AO22X1 U4622 ( .IN1(\read_value_mux[1][12] ), .IN2(n1622), .IN3(
        write_data[12]), .IN4(n3158), .Q(\words[1]/data_i[12] ) );
  AO22X1 U4623 ( .IN1(\read_value_mux[1][13] ), .IN2(n1622), .IN3(
        write_data[13]), .IN4(n3158), .Q(\words[1]/data_i[13] ) );
  AO22X1 U4624 ( .IN1(\read_value_mux[1][14] ), .IN2(n1622), .IN3(
        write_data[14]), .IN4(n3158), .Q(\words[1]/data_i[14] ) );
  AO22X1 U4625 ( .IN1(\read_value_mux[1][15] ), .IN2(n1622), .IN3(
        write_data[15]), .IN4(n3158), .Q(\words[1]/data_i[15] ) );
  AO22X1 U4626 ( .IN1(\read_value_mux[1][16] ), .IN2(n1622), .IN3(
        write_data[16]), .IN4(n3158), .Q(\words[1]/data_i[16] ) );
  AO22X1 U4627 ( .IN1(\read_value_mux[1][17] ), .IN2(n1622), .IN3(
        write_data[17]), .IN4(n3158), .Q(\words[1]/data_i[17] ) );
  AO22X1 U4628 ( .IN1(\read_value_mux[1][18] ), .IN2(n1622), .IN3(
        write_data[18]), .IN4(n3158), .Q(\words[1]/data_i[18] ) );
  AO22X1 U4629 ( .IN1(\read_value_mux[1][19] ), .IN2(n1622), .IN3(
        write_data[19]), .IN4(n3158), .Q(\words[1]/data_i[19] ) );
  AO22X1 U4630 ( .IN1(\read_value_mux[1][1] ), .IN2(n1622), .IN3(write_data[1]), .IN4(n3158), .Q(\words[1]/data_i[1] ) );
  AO22X1 U4631 ( .IN1(\read_value_mux[1][20] ), .IN2(n1622), .IN3(
        write_data[20]), .IN4(n3158), .Q(\words[1]/data_i[20] ) );
  AO22X1 U4632 ( .IN1(\read_value_mux[1][21] ), .IN2(n1622), .IN3(
        write_data[21]), .IN4(n3158), .Q(\words[1]/data_i[21] ) );
  AO22X1 U4633 ( .IN1(\read_value_mux[1][22] ), .IN2(n1622), .IN3(
        write_data[22]), .IN4(n3158), .Q(\words[1]/data_i[22] ) );
  AO22X1 U4634 ( .IN1(\read_value_mux[1][23] ), .IN2(n1622), .IN3(
        write_data[23]), .IN4(n3158), .Q(\words[1]/data_i[23] ) );
  AO22X1 U4635 ( .IN1(\read_value_mux[1][24] ), .IN2(n1622), .IN3(
        write_data[24]), .IN4(n3158), .Q(\words[1]/data_i[24] ) );
  AO22X1 U4636 ( .IN1(\read_value_mux[1][25] ), .IN2(n1622), .IN3(
        write_data[25]), .IN4(n3158), .Q(\words[1]/data_i[25] ) );
  AO22X1 U4637 ( .IN1(\read_value_mux[1][26] ), .IN2(n1622), .IN3(
        write_data[26]), .IN4(n3158), .Q(\words[1]/data_i[26] ) );
  AO22X1 U4638 ( .IN1(\read_value_mux[1][27] ), .IN2(n1622), .IN3(
        write_data[27]), .IN4(n3158), .Q(\words[1]/data_i[27] ) );
  AO22X1 U4639 ( .IN1(\read_value_mux[1][28] ), .IN2(n1622), .IN3(
        write_data[28]), .IN4(n3158), .Q(\words[1]/data_i[28] ) );
  AO22X1 U4640 ( .IN1(\read_value_mux[1][29] ), .IN2(n1622), .IN3(
        write_data[29]), .IN4(n3158), .Q(\words[1]/data_i[29] ) );
  AO22X1 U4641 ( .IN1(\read_value_mux[1][2] ), .IN2(n1622), .IN3(write_data[2]), .IN4(n3158), .Q(\words[1]/data_i[2] ) );
  AO22X1 U4642 ( .IN1(\read_value_mux[1][30] ), .IN2(n1622), .IN3(
        write_data[30]), .IN4(n3158), .Q(\words[1]/data_i[30] ) );
  AO22X1 U4643 ( .IN1(\read_value_mux[1][31] ), .IN2(n1622), .IN3(
        write_data[31]), .IN4(n3158), .Q(\words[1]/data_i[31] ) );
  AO22X1 U4644 ( .IN1(\read_value_mux[1][3] ), .IN2(n1622), .IN3(write_data[3]), .IN4(n3158), .Q(\words[1]/data_i[3] ) );
  AO22X1 U4645 ( .IN1(\read_value_mux[1][4] ), .IN2(n1622), .IN3(write_data[4]), .IN4(n3158), .Q(\words[1]/data_i[4] ) );
  AO22X1 U4646 ( .IN1(\read_value_mux[1][5] ), .IN2(n1622), .IN3(write_data[5]), .IN4(n3158), .Q(\words[1]/data_i[5] ) );
  AO22X1 U4647 ( .IN1(\read_value_mux[1][6] ), .IN2(n1622), .IN3(write_data[6]), .IN4(n3158), .Q(\words[1]/data_i[6] ) );
  AO22X1 U4648 ( .IN1(\read_value_mux[1][7] ), .IN2(n1622), .IN3(write_data[7]), .IN4(n3158), .Q(\words[1]/data_i[7] ) );
  AO22X1 U4649 ( .IN1(\read_value_mux[1][8] ), .IN2(n1622), .IN3(write_data[8]), .IN4(n3158), .Q(\words[1]/data_i[8] ) );
  AO22X1 U4650 ( .IN1(\read_value_mux[1][9] ), .IN2(n1622), .IN3(write_data[9]), .IN4(n3158), .Q(\words[1]/data_i[9] ) );
  AO21X1 U4651 ( .IN1(\words[1]/valid_o ), .IN2(n1743), .IN3(n3158), .Q(
        \words[1]/valid_i ) );
  AO22X1 U4652 ( .IN1(\read_value_mux[20][0] ), .IN2(n1628), .IN3(
        write_data[0]), .IN4(n3159), .Q(\words[20]/data_i[0] ) );
  AO22X1 U4653 ( .IN1(\read_value_mux[20][10] ), .IN2(n1628), .IN3(
        write_data[10]), .IN4(n3159), .Q(\words[20]/data_i[10] ) );
  AO22X1 U4654 ( .IN1(\read_value_mux[20][11] ), .IN2(n1628), .IN3(
        write_data[11]), .IN4(n3159), .Q(\words[20]/data_i[11] ) );
  AO22X1 U4655 ( .IN1(\read_value_mux[20][12] ), .IN2(n1628), .IN3(
        write_data[12]), .IN4(n3159), .Q(\words[20]/data_i[12] ) );
  AO22X1 U4656 ( .IN1(\read_value_mux[20][13] ), .IN2(n1628), .IN3(
        write_data[13]), .IN4(n3159), .Q(\words[20]/data_i[13] ) );
  AO22X1 U4657 ( .IN1(\read_value_mux[20][14] ), .IN2(n1628), .IN3(
        write_data[14]), .IN4(n3159), .Q(\words[20]/data_i[14] ) );
  AO22X1 U4658 ( .IN1(\read_value_mux[20][15] ), .IN2(n1628), .IN3(
        write_data[15]), .IN4(n3159), .Q(\words[20]/data_i[15] ) );
  AO22X1 U4659 ( .IN1(\read_value_mux[20][16] ), .IN2(n1628), .IN3(
        write_data[16]), .IN4(n3159), .Q(\words[20]/data_i[16] ) );
  AO22X1 U4660 ( .IN1(\read_value_mux[20][17] ), .IN2(n1628), .IN3(
        write_data[17]), .IN4(n3159), .Q(\words[20]/data_i[17] ) );
  AO22X1 U4661 ( .IN1(\read_value_mux[20][18] ), .IN2(n1628), .IN3(
        write_data[18]), .IN4(n3159), .Q(\words[20]/data_i[18] ) );
  AO22X1 U4662 ( .IN1(\read_value_mux[20][19] ), .IN2(n1628), .IN3(
        write_data[19]), .IN4(n3159), .Q(\words[20]/data_i[19] ) );
  AO22X1 U4663 ( .IN1(\read_value_mux[20][1] ), .IN2(n1628), .IN3(
        write_data[1]), .IN4(n3159), .Q(\words[20]/data_i[1] ) );
  AO22X1 U4664 ( .IN1(\read_value_mux[20][20] ), .IN2(n1628), .IN3(
        write_data[20]), .IN4(n3159), .Q(\words[20]/data_i[20] ) );
  AO22X1 U4665 ( .IN1(\read_value_mux[20][21] ), .IN2(n1628), .IN3(
        write_data[21]), .IN4(n3159), .Q(\words[20]/data_i[21] ) );
  AO22X1 U4666 ( .IN1(\read_value_mux[20][22] ), .IN2(n1628), .IN3(
        write_data[22]), .IN4(n3159), .Q(\words[20]/data_i[22] ) );
  AO22X1 U4667 ( .IN1(\read_value_mux[20][23] ), .IN2(n1628), .IN3(
        write_data[23]), .IN4(n3159), .Q(\words[20]/data_i[23] ) );
  AO22X1 U4668 ( .IN1(\read_value_mux[20][24] ), .IN2(n1628), .IN3(
        write_data[24]), .IN4(n3159), .Q(\words[20]/data_i[24] ) );
  AO22X1 U4669 ( .IN1(\read_value_mux[20][25] ), .IN2(n1628), .IN3(
        write_data[25]), .IN4(n3159), .Q(\words[20]/data_i[25] ) );
  AO22X1 U4670 ( .IN1(\read_value_mux[20][26] ), .IN2(n1628), .IN3(
        write_data[26]), .IN4(n3159), .Q(\words[20]/data_i[26] ) );
  AO22X1 U4671 ( .IN1(\read_value_mux[20][27] ), .IN2(n1628), .IN3(
        write_data[27]), .IN4(n3159), .Q(\words[20]/data_i[27] ) );
  AO22X1 U4672 ( .IN1(\read_value_mux[20][28] ), .IN2(n1628), .IN3(
        write_data[28]), .IN4(n3159), .Q(\words[20]/data_i[28] ) );
  AO22X1 U4673 ( .IN1(\read_value_mux[20][29] ), .IN2(n1628), .IN3(
        write_data[29]), .IN4(n3159), .Q(\words[20]/data_i[29] ) );
  AO22X1 U4674 ( .IN1(\read_value_mux[20][2] ), .IN2(n1628), .IN3(
        write_data[2]), .IN4(n3159), .Q(\words[20]/data_i[2] ) );
  AO22X1 U4675 ( .IN1(\read_value_mux[20][30] ), .IN2(n1628), .IN3(
        write_data[30]), .IN4(n3159), .Q(\words[20]/data_i[30] ) );
  AO22X1 U4676 ( .IN1(\read_value_mux[20][31] ), .IN2(n1628), .IN3(
        write_data[31]), .IN4(n3159), .Q(\words[20]/data_i[31] ) );
  AO22X1 U4677 ( .IN1(\read_value_mux[20][3] ), .IN2(n1628), .IN3(
        write_data[3]), .IN4(n3159), .Q(\words[20]/data_i[3] ) );
  AO22X1 U4678 ( .IN1(\read_value_mux[20][4] ), .IN2(n1628), .IN3(
        write_data[4]), .IN4(n3159), .Q(\words[20]/data_i[4] ) );
  AO22X1 U4679 ( .IN1(\read_value_mux[20][5] ), .IN2(n1628), .IN3(
        write_data[5]), .IN4(n3159), .Q(\words[20]/data_i[5] ) );
  AO22X1 U4680 ( .IN1(\read_value_mux[20][6] ), .IN2(n1628), .IN3(
        write_data[6]), .IN4(n3159), .Q(\words[20]/data_i[6] ) );
  AO22X1 U4681 ( .IN1(\read_value_mux[20][7] ), .IN2(n1628), .IN3(
        write_data[7]), .IN4(n3159), .Q(\words[20]/data_i[7] ) );
  AO22X1 U4682 ( .IN1(\read_value_mux[20][8] ), .IN2(n1628), .IN3(
        write_data[8]), .IN4(n3159), .Q(\words[20]/data_i[8] ) );
  AO22X1 U4683 ( .IN1(\read_value_mux[20][9] ), .IN2(n1628), .IN3(
        write_data[9]), .IN4(n3159), .Q(\words[20]/data_i[9] ) );
  AO21X1 U4684 ( .IN1(\words[20]/valid_o ), .IN2(n1743), .IN3(n3159), .Q(
        \words[20]/valid_i ) );
  AO22X1 U4685 ( .IN1(\read_value_mux[21][0] ), .IN2(n1629), .IN3(
        write_data[0]), .IN4(n3160), .Q(\words[21]/data_i[0] ) );
  AO22X1 U4686 ( .IN1(\read_value_mux[21][10] ), .IN2(n1629), .IN3(
        write_data[10]), .IN4(n3160), .Q(\words[21]/data_i[10] ) );
  AO22X1 U4687 ( .IN1(\read_value_mux[21][11] ), .IN2(n1629), .IN3(
        write_data[11]), .IN4(n3160), .Q(\words[21]/data_i[11] ) );
  AO22X1 U4688 ( .IN1(\read_value_mux[21][12] ), .IN2(n1629), .IN3(
        write_data[12]), .IN4(n3160), .Q(\words[21]/data_i[12] ) );
  AO22X1 U4689 ( .IN1(\read_value_mux[21][13] ), .IN2(n1629), .IN3(
        write_data[13]), .IN4(n3160), .Q(\words[21]/data_i[13] ) );
  AO22X1 U4690 ( .IN1(\read_value_mux[21][14] ), .IN2(n1629), .IN3(
        write_data[14]), .IN4(n3160), .Q(\words[21]/data_i[14] ) );
  AO22X1 U4691 ( .IN1(\read_value_mux[21][15] ), .IN2(n1629), .IN3(
        write_data[15]), .IN4(n3160), .Q(\words[21]/data_i[15] ) );
  AO22X1 U4692 ( .IN1(\read_value_mux[21][16] ), .IN2(n1629), .IN3(
        write_data[16]), .IN4(n3160), .Q(\words[21]/data_i[16] ) );
  AO22X1 U4693 ( .IN1(\read_value_mux[21][17] ), .IN2(n1629), .IN3(
        write_data[17]), .IN4(n3160), .Q(\words[21]/data_i[17] ) );
  AO22X1 U4694 ( .IN1(\read_value_mux[21][18] ), .IN2(n1629), .IN3(
        write_data[18]), .IN4(n3160), .Q(\words[21]/data_i[18] ) );
  AO22X1 U4695 ( .IN1(\read_value_mux[21][19] ), .IN2(n1629), .IN3(
        write_data[19]), .IN4(n3160), .Q(\words[21]/data_i[19] ) );
  AO22X1 U4696 ( .IN1(\read_value_mux[21][1] ), .IN2(n1629), .IN3(
        write_data[1]), .IN4(n3160), .Q(\words[21]/data_i[1] ) );
  AO22X1 U4697 ( .IN1(\read_value_mux[21][20] ), .IN2(n1629), .IN3(
        write_data[20]), .IN4(n3160), .Q(\words[21]/data_i[20] ) );
  AO22X1 U4698 ( .IN1(\read_value_mux[21][21] ), .IN2(n1629), .IN3(
        write_data[21]), .IN4(n3160), .Q(\words[21]/data_i[21] ) );
  AO22X1 U4699 ( .IN1(\read_value_mux[21][22] ), .IN2(n1629), .IN3(
        write_data[22]), .IN4(n3160), .Q(\words[21]/data_i[22] ) );
  AO22X1 U4700 ( .IN1(\read_value_mux[21][23] ), .IN2(n1629), .IN3(
        write_data[23]), .IN4(n3160), .Q(\words[21]/data_i[23] ) );
  AO22X1 U4701 ( .IN1(\read_value_mux[21][24] ), .IN2(n1629), .IN3(
        write_data[24]), .IN4(n3160), .Q(\words[21]/data_i[24] ) );
  AO22X1 U4702 ( .IN1(\read_value_mux[21][25] ), .IN2(n1629), .IN3(
        write_data[25]), .IN4(n3160), .Q(\words[21]/data_i[25] ) );
  AO22X1 U4703 ( .IN1(\read_value_mux[21][26] ), .IN2(n1629), .IN3(
        write_data[26]), .IN4(n3160), .Q(\words[21]/data_i[26] ) );
  AO22X1 U4704 ( .IN1(\read_value_mux[21][27] ), .IN2(n1629), .IN3(
        write_data[27]), .IN4(n3160), .Q(\words[21]/data_i[27] ) );
  AO22X1 U4705 ( .IN1(\read_value_mux[21][28] ), .IN2(n1629), .IN3(
        write_data[28]), .IN4(n3160), .Q(\words[21]/data_i[28] ) );
  AO22X1 U4706 ( .IN1(\read_value_mux[21][29] ), .IN2(n1629), .IN3(
        write_data[29]), .IN4(n3160), .Q(\words[21]/data_i[29] ) );
  AO22X1 U4707 ( .IN1(\read_value_mux[21][2] ), .IN2(n1629), .IN3(
        write_data[2]), .IN4(n3160), .Q(\words[21]/data_i[2] ) );
  AO22X1 U4708 ( .IN1(\read_value_mux[21][30] ), .IN2(n1629), .IN3(
        write_data[30]), .IN4(n3160), .Q(\words[21]/data_i[30] ) );
  AO22X1 U4709 ( .IN1(\read_value_mux[21][31] ), .IN2(n1629), .IN3(
        write_data[31]), .IN4(n3160), .Q(\words[21]/data_i[31] ) );
  AO22X1 U4710 ( .IN1(\read_value_mux[21][3] ), .IN2(n1629), .IN3(
        write_data[3]), .IN4(n3160), .Q(\words[21]/data_i[3] ) );
  AO22X1 U4711 ( .IN1(\read_value_mux[21][4] ), .IN2(n1629), .IN3(
        write_data[4]), .IN4(n3160), .Q(\words[21]/data_i[4] ) );
  AO22X1 U4712 ( .IN1(\read_value_mux[21][5] ), .IN2(n1629), .IN3(
        write_data[5]), .IN4(n3160), .Q(\words[21]/data_i[5] ) );
  AO22X1 U4713 ( .IN1(\read_value_mux[21][6] ), .IN2(n1629), .IN3(
        write_data[6]), .IN4(n3160), .Q(\words[21]/data_i[6] ) );
  AO22X1 U4714 ( .IN1(\read_value_mux[21][7] ), .IN2(n1629), .IN3(
        write_data[7]), .IN4(n3160), .Q(\words[21]/data_i[7] ) );
  AO22X1 U4715 ( .IN1(\read_value_mux[21][8] ), .IN2(n1629), .IN3(
        write_data[8]), .IN4(n3160), .Q(\words[21]/data_i[8] ) );
  AO22X1 U4716 ( .IN1(\read_value_mux[21][9] ), .IN2(n1629), .IN3(
        write_data[9]), .IN4(n3160), .Q(\words[21]/data_i[9] ) );
  AO21X1 U4717 ( .IN1(\words[21]/valid_o ), .IN2(n1743), .IN3(n3160), .Q(
        \words[21]/valid_i ) );
  AO22X1 U4718 ( .IN1(\read_value_mux[22][0] ), .IN2(n1637), .IN3(
        write_data[0]), .IN4(n3161), .Q(\words[22]/data_i[0] ) );
  AO22X1 U4719 ( .IN1(\read_value_mux[22][10] ), .IN2(n1637), .IN3(
        write_data[10]), .IN4(n3161), .Q(\words[22]/data_i[10] ) );
  AO22X1 U4720 ( .IN1(\read_value_mux[22][11] ), .IN2(n1637), .IN3(
        write_data[11]), .IN4(n3161), .Q(\words[22]/data_i[11] ) );
  AO22X1 U4721 ( .IN1(\read_value_mux[22][12] ), .IN2(n1637), .IN3(
        write_data[12]), .IN4(n3161), .Q(\words[22]/data_i[12] ) );
  AO22X1 U4722 ( .IN1(\read_value_mux[22][13] ), .IN2(n1637), .IN3(
        write_data[13]), .IN4(n3161), .Q(\words[22]/data_i[13] ) );
  AO22X1 U4723 ( .IN1(\read_value_mux[22][14] ), .IN2(n1637), .IN3(
        write_data[14]), .IN4(n3161), .Q(\words[22]/data_i[14] ) );
  AO22X1 U4724 ( .IN1(\read_value_mux[22][15] ), .IN2(n1637), .IN3(
        write_data[15]), .IN4(n3161), .Q(\words[22]/data_i[15] ) );
  AO22X1 U4725 ( .IN1(\read_value_mux[22][16] ), .IN2(n1637), .IN3(
        write_data[16]), .IN4(n3161), .Q(\words[22]/data_i[16] ) );
  AO22X1 U4726 ( .IN1(\read_value_mux[22][17] ), .IN2(n1637), .IN3(
        write_data[17]), .IN4(n3161), .Q(\words[22]/data_i[17] ) );
  AO22X1 U4727 ( .IN1(\read_value_mux[22][18] ), .IN2(n1637), .IN3(
        write_data[18]), .IN4(n3161), .Q(\words[22]/data_i[18] ) );
  AO22X1 U4728 ( .IN1(\read_value_mux[22][19] ), .IN2(n1637), .IN3(
        write_data[19]), .IN4(n3161), .Q(\words[22]/data_i[19] ) );
  AO22X1 U4729 ( .IN1(\read_value_mux[22][1] ), .IN2(n1637), .IN3(
        write_data[1]), .IN4(n3161), .Q(\words[22]/data_i[1] ) );
  AO22X1 U4730 ( .IN1(\read_value_mux[22][20] ), .IN2(n1637), .IN3(
        write_data[20]), .IN4(n3161), .Q(\words[22]/data_i[20] ) );
  AO22X1 U4731 ( .IN1(\read_value_mux[22][21] ), .IN2(n1637), .IN3(
        write_data[21]), .IN4(n3161), .Q(\words[22]/data_i[21] ) );
  AO22X1 U4732 ( .IN1(\read_value_mux[22][22] ), .IN2(n1637), .IN3(
        write_data[22]), .IN4(n3161), .Q(\words[22]/data_i[22] ) );
  AO22X1 U4733 ( .IN1(\read_value_mux[22][23] ), .IN2(n1637), .IN3(
        write_data[23]), .IN4(n3161), .Q(\words[22]/data_i[23] ) );
  AO22X1 U4734 ( .IN1(\read_value_mux[22][24] ), .IN2(n1637), .IN3(
        write_data[24]), .IN4(n3161), .Q(\words[22]/data_i[24] ) );
  AO22X1 U4735 ( .IN1(\read_value_mux[22][25] ), .IN2(n1637), .IN3(
        write_data[25]), .IN4(n3161), .Q(\words[22]/data_i[25] ) );
  AO22X1 U4736 ( .IN1(\read_value_mux[22][26] ), .IN2(n1637), .IN3(
        write_data[26]), .IN4(n3161), .Q(\words[22]/data_i[26] ) );
  AO22X1 U4737 ( .IN1(\read_value_mux[22][27] ), .IN2(n1637), .IN3(
        write_data[27]), .IN4(n3161), .Q(\words[22]/data_i[27] ) );
  AO22X1 U4738 ( .IN1(\read_value_mux[22][28] ), .IN2(n1637), .IN3(
        write_data[28]), .IN4(n3161), .Q(\words[22]/data_i[28] ) );
  AO22X1 U4739 ( .IN1(\read_value_mux[22][29] ), .IN2(n1637), .IN3(
        write_data[29]), .IN4(n3161), .Q(\words[22]/data_i[29] ) );
  AO22X1 U4740 ( .IN1(\read_value_mux[22][2] ), .IN2(n1637), .IN3(
        write_data[2]), .IN4(n3161), .Q(\words[22]/data_i[2] ) );
  AO22X1 U4741 ( .IN1(\read_value_mux[22][30] ), .IN2(n1637), .IN3(
        write_data[30]), .IN4(n3161), .Q(\words[22]/data_i[30] ) );
  AO22X1 U4742 ( .IN1(\read_value_mux[22][31] ), .IN2(n1637), .IN3(
        write_data[31]), .IN4(n3161), .Q(\words[22]/data_i[31] ) );
  AO22X1 U4743 ( .IN1(\read_value_mux[22][3] ), .IN2(n1637), .IN3(
        write_data[3]), .IN4(n3161), .Q(\words[22]/data_i[3] ) );
  AO22X1 U4744 ( .IN1(\read_value_mux[22][4] ), .IN2(n1637), .IN3(
        write_data[4]), .IN4(n3161), .Q(\words[22]/data_i[4] ) );
  AO22X1 U4745 ( .IN1(\read_value_mux[22][5] ), .IN2(n1637), .IN3(
        write_data[5]), .IN4(n3161), .Q(\words[22]/data_i[5] ) );
  AO22X1 U4746 ( .IN1(\read_value_mux[22][6] ), .IN2(n1637), .IN3(
        write_data[6]), .IN4(n3161), .Q(\words[22]/data_i[6] ) );
  AO22X1 U4747 ( .IN1(\read_value_mux[22][7] ), .IN2(n1637), .IN3(
        write_data[7]), .IN4(n3161), .Q(\words[22]/data_i[7] ) );
  AO22X1 U4748 ( .IN1(\read_value_mux[22][8] ), .IN2(n1637), .IN3(
        write_data[8]), .IN4(n3161), .Q(\words[22]/data_i[8] ) );
  AO22X1 U4749 ( .IN1(\read_value_mux[22][9] ), .IN2(n1637), .IN3(
        write_data[9]), .IN4(n3161), .Q(\words[22]/data_i[9] ) );
  AO21X1 U4750 ( .IN1(\words[22]/valid_o ), .IN2(n1743), .IN3(n3161), .Q(
        \words[22]/valid_i ) );
  AO22X1 U4751 ( .IN1(\read_value_mux[23][0] ), .IN2(n1638), .IN3(
        write_data[0]), .IN4(n3163), .Q(\words[23]/data_i[0] ) );
  AO22X1 U4752 ( .IN1(\read_value_mux[23][10] ), .IN2(n1638), .IN3(
        write_data[10]), .IN4(n3163), .Q(\words[23]/data_i[10] ) );
  AO22X1 U4753 ( .IN1(\read_value_mux[23][11] ), .IN2(n1638), .IN3(
        write_data[11]), .IN4(n3163), .Q(\words[23]/data_i[11] ) );
  AO22X1 U4754 ( .IN1(\read_value_mux[23][12] ), .IN2(n1638), .IN3(
        write_data[12]), .IN4(n3163), .Q(\words[23]/data_i[12] ) );
  AO22X1 U4755 ( .IN1(\read_value_mux[23][13] ), .IN2(n1638), .IN3(
        write_data[13]), .IN4(n3163), .Q(\words[23]/data_i[13] ) );
  AO22X1 U4756 ( .IN1(\read_value_mux[23][14] ), .IN2(n1638), .IN3(
        write_data[14]), .IN4(n3163), .Q(\words[23]/data_i[14] ) );
  AO22X1 U4757 ( .IN1(\read_value_mux[23][15] ), .IN2(n1638), .IN3(
        write_data[15]), .IN4(n3163), .Q(\words[23]/data_i[15] ) );
  AO22X1 U4758 ( .IN1(\read_value_mux[23][16] ), .IN2(n1638), .IN3(
        write_data[16]), .IN4(n3163), .Q(\words[23]/data_i[16] ) );
  AO22X1 U4759 ( .IN1(\read_value_mux[23][17] ), .IN2(n1638), .IN3(
        write_data[17]), .IN4(n3163), .Q(\words[23]/data_i[17] ) );
  AO22X1 U4760 ( .IN1(\read_value_mux[23][18] ), .IN2(n1638), .IN3(
        write_data[18]), .IN4(n3163), .Q(\words[23]/data_i[18] ) );
  AO22X1 U4761 ( .IN1(\read_value_mux[23][19] ), .IN2(n1638), .IN3(
        write_data[19]), .IN4(n3163), .Q(\words[23]/data_i[19] ) );
  AO22X1 U4762 ( .IN1(\read_value_mux[23][1] ), .IN2(n1638), .IN3(
        write_data[1]), .IN4(n3163), .Q(\words[23]/data_i[1] ) );
  AO22X1 U4763 ( .IN1(\read_value_mux[23][20] ), .IN2(n1638), .IN3(
        write_data[20]), .IN4(n3163), .Q(\words[23]/data_i[20] ) );
  AO22X1 U4764 ( .IN1(\read_value_mux[23][21] ), .IN2(n1638), .IN3(
        write_data[21]), .IN4(n3163), .Q(\words[23]/data_i[21] ) );
  AO22X1 U4765 ( .IN1(\read_value_mux[23][22] ), .IN2(n1638), .IN3(
        write_data[22]), .IN4(n3163), .Q(\words[23]/data_i[22] ) );
  AO22X1 U4766 ( .IN1(\read_value_mux[23][23] ), .IN2(n1638), .IN3(
        write_data[23]), .IN4(n3163), .Q(\words[23]/data_i[23] ) );
  AO22X1 U4767 ( .IN1(\read_value_mux[23][24] ), .IN2(n1638), .IN3(
        write_data[24]), .IN4(n3163), .Q(\words[23]/data_i[24] ) );
  AO22X1 U4768 ( .IN1(\read_value_mux[23][25] ), .IN2(n1638), .IN3(
        write_data[25]), .IN4(n3163), .Q(\words[23]/data_i[25] ) );
  AO22X1 U4769 ( .IN1(\read_value_mux[23][26] ), .IN2(n1638), .IN3(
        write_data[26]), .IN4(n3163), .Q(\words[23]/data_i[26] ) );
  AO22X1 U4770 ( .IN1(\read_value_mux[23][27] ), .IN2(n1638), .IN3(
        write_data[27]), .IN4(n3163), .Q(\words[23]/data_i[27] ) );
  AO22X1 U4771 ( .IN1(\read_value_mux[23][28] ), .IN2(n1638), .IN3(
        write_data[28]), .IN4(n3163), .Q(\words[23]/data_i[28] ) );
  AO22X1 U4772 ( .IN1(\read_value_mux[23][29] ), .IN2(n1638), .IN3(
        write_data[29]), .IN4(n3163), .Q(\words[23]/data_i[29] ) );
  AO22X1 U4773 ( .IN1(\read_value_mux[23][2] ), .IN2(n1638), .IN3(
        write_data[2]), .IN4(n3163), .Q(\words[23]/data_i[2] ) );
  AO22X1 U4774 ( .IN1(\read_value_mux[23][30] ), .IN2(n1638), .IN3(
        write_data[30]), .IN4(n3163), .Q(\words[23]/data_i[30] ) );
  AO22X1 U4775 ( .IN1(\read_value_mux[23][31] ), .IN2(n1638), .IN3(
        write_data[31]), .IN4(n3163), .Q(\words[23]/data_i[31] ) );
  AO22X1 U4776 ( .IN1(\read_value_mux[23][3] ), .IN2(n1638), .IN3(
        write_data[3]), .IN4(n3163), .Q(\words[23]/data_i[3] ) );
  AO22X1 U4777 ( .IN1(\read_value_mux[23][4] ), .IN2(n1638), .IN3(
        write_data[4]), .IN4(n3163), .Q(\words[23]/data_i[4] ) );
  AO22X1 U4778 ( .IN1(\read_value_mux[23][5] ), .IN2(n1638), .IN3(
        write_data[5]), .IN4(n3163), .Q(\words[23]/data_i[5] ) );
  AO22X1 U4779 ( .IN1(\read_value_mux[23][6] ), .IN2(n1638), .IN3(
        write_data[6]), .IN4(n3163), .Q(\words[23]/data_i[6] ) );
  AO22X1 U4780 ( .IN1(\read_value_mux[23][7] ), .IN2(n1638), .IN3(
        write_data[7]), .IN4(n3163), .Q(\words[23]/data_i[7] ) );
  AO22X1 U4781 ( .IN1(\read_value_mux[23][8] ), .IN2(n1638), .IN3(
        write_data[8]), .IN4(n3163), .Q(\words[23]/data_i[8] ) );
  AO22X1 U4782 ( .IN1(\read_value_mux[23][9] ), .IN2(n1638), .IN3(
        write_data[9]), .IN4(n3163), .Q(\words[23]/data_i[9] ) );
  AO21X1 U4783 ( .IN1(\words[23]/valid_o ), .IN2(n1743), .IN3(n3163), .Q(
        \words[23]/valid_i ) );
  AO22X1 U4784 ( .IN1(\read_value_mux[24][0] ), .IN2(n1630), .IN3(
        write_data[0]), .IN4(n3165), .Q(\words[24]/data_i[0] ) );
  AO22X1 U4785 ( .IN1(\read_value_mux[24][10] ), .IN2(n1630), .IN3(
        write_data[10]), .IN4(n3165), .Q(\words[24]/data_i[10] ) );
  AO22X1 U4786 ( .IN1(\read_value_mux[24][11] ), .IN2(n1630), .IN3(
        write_data[11]), .IN4(n3165), .Q(\words[24]/data_i[11] ) );
  AO22X1 U4787 ( .IN1(\read_value_mux[24][12] ), .IN2(n1630), .IN3(
        write_data[12]), .IN4(n3165), .Q(\words[24]/data_i[12] ) );
  AO22X1 U4788 ( .IN1(\read_value_mux[24][13] ), .IN2(n1630), .IN3(
        write_data[13]), .IN4(n3165), .Q(\words[24]/data_i[13] ) );
  AO22X1 U4789 ( .IN1(\read_value_mux[24][14] ), .IN2(n1630), .IN3(
        write_data[14]), .IN4(n3165), .Q(\words[24]/data_i[14] ) );
  AO22X1 U4790 ( .IN1(\read_value_mux[24][15] ), .IN2(n1630), .IN3(
        write_data[15]), .IN4(n3165), .Q(\words[24]/data_i[15] ) );
  AO22X1 U4791 ( .IN1(\read_value_mux[24][16] ), .IN2(n1630), .IN3(
        write_data[16]), .IN4(n3165), .Q(\words[24]/data_i[16] ) );
  AO22X1 U4792 ( .IN1(\read_value_mux[24][17] ), .IN2(n1630), .IN3(
        write_data[17]), .IN4(n3165), .Q(\words[24]/data_i[17] ) );
  AO22X1 U4793 ( .IN1(\read_value_mux[24][18] ), .IN2(n1630), .IN3(
        write_data[18]), .IN4(n3165), .Q(\words[24]/data_i[18] ) );
  AO22X1 U4794 ( .IN1(\read_value_mux[24][19] ), .IN2(n1630), .IN3(
        write_data[19]), .IN4(n3165), .Q(\words[24]/data_i[19] ) );
  AO22X1 U4795 ( .IN1(\read_value_mux[24][1] ), .IN2(n1630), .IN3(
        write_data[1]), .IN4(n3165), .Q(\words[24]/data_i[1] ) );
  AO22X1 U4796 ( .IN1(\read_value_mux[24][20] ), .IN2(n1630), .IN3(
        write_data[20]), .IN4(n3165), .Q(\words[24]/data_i[20] ) );
  AO22X1 U4797 ( .IN1(\read_value_mux[24][21] ), .IN2(n1630), .IN3(
        write_data[21]), .IN4(n3165), .Q(\words[24]/data_i[21] ) );
  AO22X1 U4798 ( .IN1(\read_value_mux[24][22] ), .IN2(n1630), .IN3(
        write_data[22]), .IN4(n3165), .Q(\words[24]/data_i[22] ) );
  AO22X1 U4799 ( .IN1(\read_value_mux[24][23] ), .IN2(n1630), .IN3(
        write_data[23]), .IN4(n3165), .Q(\words[24]/data_i[23] ) );
  AO22X1 U4800 ( .IN1(\read_value_mux[24][24] ), .IN2(n1630), .IN3(
        write_data[24]), .IN4(n3165), .Q(\words[24]/data_i[24] ) );
  AO22X1 U4801 ( .IN1(\read_value_mux[24][25] ), .IN2(n1630), .IN3(
        write_data[25]), .IN4(n3165), .Q(\words[24]/data_i[25] ) );
  AO22X1 U4802 ( .IN1(\read_value_mux[24][26] ), .IN2(n1630), .IN3(
        write_data[26]), .IN4(n3165), .Q(\words[24]/data_i[26] ) );
  AO22X1 U4803 ( .IN1(\read_value_mux[24][27] ), .IN2(n1630), .IN3(
        write_data[27]), .IN4(n3165), .Q(\words[24]/data_i[27] ) );
  AO22X1 U4804 ( .IN1(\read_value_mux[24][28] ), .IN2(n1630), .IN3(
        write_data[28]), .IN4(n3165), .Q(\words[24]/data_i[28] ) );
  AO22X1 U4805 ( .IN1(\read_value_mux[24][29] ), .IN2(n1630), .IN3(
        write_data[29]), .IN4(n3165), .Q(\words[24]/data_i[29] ) );
  AO22X1 U4806 ( .IN1(\read_value_mux[24][2] ), .IN2(n1630), .IN3(
        write_data[2]), .IN4(n3165), .Q(\words[24]/data_i[2] ) );
  AO22X1 U4807 ( .IN1(\read_value_mux[24][30] ), .IN2(n1630), .IN3(
        write_data[30]), .IN4(n3165), .Q(\words[24]/data_i[30] ) );
  AO22X1 U4808 ( .IN1(\read_value_mux[24][31] ), .IN2(n1630), .IN3(
        write_data[31]), .IN4(n3165), .Q(\words[24]/data_i[31] ) );
  AO22X1 U4809 ( .IN1(\read_value_mux[24][3] ), .IN2(n1630), .IN3(
        write_data[3]), .IN4(n3165), .Q(\words[24]/data_i[3] ) );
  AO22X1 U4810 ( .IN1(\read_value_mux[24][4] ), .IN2(n1630), .IN3(
        write_data[4]), .IN4(n3165), .Q(\words[24]/data_i[4] ) );
  AO22X1 U4811 ( .IN1(\read_value_mux[24][5] ), .IN2(n1630), .IN3(
        write_data[5]), .IN4(n3165), .Q(\words[24]/data_i[5] ) );
  AO22X1 U4812 ( .IN1(\read_value_mux[24][6] ), .IN2(n1630), .IN3(
        write_data[6]), .IN4(n3165), .Q(\words[24]/data_i[6] ) );
  AO22X1 U4813 ( .IN1(\read_value_mux[24][7] ), .IN2(n1630), .IN3(
        write_data[7]), .IN4(n3165), .Q(\words[24]/data_i[7] ) );
  AO22X1 U4814 ( .IN1(\read_value_mux[24][8] ), .IN2(n1630), .IN3(
        write_data[8]), .IN4(n3165), .Q(\words[24]/data_i[8] ) );
  AO22X1 U4815 ( .IN1(\read_value_mux[24][9] ), .IN2(n1630), .IN3(
        write_data[9]), .IN4(n3165), .Q(\words[24]/data_i[9] ) );
  AO21X1 U4816 ( .IN1(\words[24]/valid_o ), .IN2(n1743), .IN3(n3165), .Q(
        \words[24]/valid_i ) );
  AO22X1 U4817 ( .IN1(\read_value_mux[25][0] ), .IN2(n1631), .IN3(
        write_data[0]), .IN4(n3166), .Q(\words[25]/data_i[0] ) );
  AO22X1 U4818 ( .IN1(\read_value_mux[25][10] ), .IN2(n1631), .IN3(
        write_data[10]), .IN4(n3166), .Q(\words[25]/data_i[10] ) );
  AO22X1 U4819 ( .IN1(\read_value_mux[25][11] ), .IN2(n1631), .IN3(
        write_data[11]), .IN4(n3166), .Q(\words[25]/data_i[11] ) );
  AO22X1 U4820 ( .IN1(\read_value_mux[25][12] ), .IN2(n1631), .IN3(
        write_data[12]), .IN4(n3166), .Q(\words[25]/data_i[12] ) );
  AO22X1 U4821 ( .IN1(\read_value_mux[25][13] ), .IN2(n1631), .IN3(
        write_data[13]), .IN4(n3166), .Q(\words[25]/data_i[13] ) );
  AO22X1 U4822 ( .IN1(\read_value_mux[25][14] ), .IN2(n1631), .IN3(
        write_data[14]), .IN4(n3166), .Q(\words[25]/data_i[14] ) );
  AO22X1 U4823 ( .IN1(\read_value_mux[25][15] ), .IN2(n1631), .IN3(
        write_data[15]), .IN4(n3166), .Q(\words[25]/data_i[15] ) );
  AO22X1 U4824 ( .IN1(\read_value_mux[25][16] ), .IN2(n1631), .IN3(
        write_data[16]), .IN4(n3166), .Q(\words[25]/data_i[16] ) );
  AO22X1 U4825 ( .IN1(\read_value_mux[25][17] ), .IN2(n1631), .IN3(
        write_data[17]), .IN4(n3166), .Q(\words[25]/data_i[17] ) );
  AO22X1 U4826 ( .IN1(\read_value_mux[25][18] ), .IN2(n1631), .IN3(
        write_data[18]), .IN4(n3166), .Q(\words[25]/data_i[18] ) );
  AO22X1 U4827 ( .IN1(\read_value_mux[25][19] ), .IN2(n1631), .IN3(
        write_data[19]), .IN4(n3166), .Q(\words[25]/data_i[19] ) );
  AO22X1 U4828 ( .IN1(\read_value_mux[25][1] ), .IN2(n1631), .IN3(
        write_data[1]), .IN4(n3166), .Q(\words[25]/data_i[1] ) );
  AO22X1 U4829 ( .IN1(\read_value_mux[25][20] ), .IN2(n1631), .IN3(
        write_data[20]), .IN4(n3166), .Q(\words[25]/data_i[20] ) );
  AO22X1 U4830 ( .IN1(\read_value_mux[25][21] ), .IN2(n1631), .IN3(
        write_data[21]), .IN4(n3166), .Q(\words[25]/data_i[21] ) );
  AO22X1 U4831 ( .IN1(\read_value_mux[25][22] ), .IN2(n1631), .IN3(
        write_data[22]), .IN4(n3166), .Q(\words[25]/data_i[22] ) );
  AO22X1 U4832 ( .IN1(\read_value_mux[25][23] ), .IN2(n1631), .IN3(
        write_data[23]), .IN4(n3166), .Q(\words[25]/data_i[23] ) );
  AO22X1 U4833 ( .IN1(\read_value_mux[25][24] ), .IN2(n1631), .IN3(
        write_data[24]), .IN4(n3166), .Q(\words[25]/data_i[24] ) );
  AO22X1 U4834 ( .IN1(\read_value_mux[25][25] ), .IN2(n1631), .IN3(
        write_data[25]), .IN4(n3166), .Q(\words[25]/data_i[25] ) );
  AO22X1 U4835 ( .IN1(\read_value_mux[25][26] ), .IN2(n1631), .IN3(
        write_data[26]), .IN4(n3166), .Q(\words[25]/data_i[26] ) );
  AO22X1 U4836 ( .IN1(\read_value_mux[25][27] ), .IN2(n1631), .IN3(
        write_data[27]), .IN4(n3166), .Q(\words[25]/data_i[27] ) );
  AO22X1 U4837 ( .IN1(\read_value_mux[25][28] ), .IN2(n1631), .IN3(
        write_data[28]), .IN4(n3166), .Q(\words[25]/data_i[28] ) );
  AO22X1 U4838 ( .IN1(\read_value_mux[25][29] ), .IN2(n1631), .IN3(
        write_data[29]), .IN4(n3166), .Q(\words[25]/data_i[29] ) );
  AO22X1 U4839 ( .IN1(\read_value_mux[25][2] ), .IN2(n1631), .IN3(
        write_data[2]), .IN4(n3166), .Q(\words[25]/data_i[2] ) );
  AO22X1 U4840 ( .IN1(\read_value_mux[25][30] ), .IN2(n1631), .IN3(
        write_data[30]), .IN4(n3166), .Q(\words[25]/data_i[30] ) );
  AO22X1 U4841 ( .IN1(\read_value_mux[25][31] ), .IN2(n1631), .IN3(
        write_data[31]), .IN4(n3166), .Q(\words[25]/data_i[31] ) );
  AO22X1 U4842 ( .IN1(\read_value_mux[25][3] ), .IN2(n1631), .IN3(
        write_data[3]), .IN4(n3166), .Q(\words[25]/data_i[3] ) );
  AO22X1 U4843 ( .IN1(\read_value_mux[25][4] ), .IN2(n1631), .IN3(
        write_data[4]), .IN4(n3166), .Q(\words[25]/data_i[4] ) );
  AO22X1 U4844 ( .IN1(\read_value_mux[25][5] ), .IN2(n1631), .IN3(
        write_data[5]), .IN4(n3166), .Q(\words[25]/data_i[5] ) );
  AO22X1 U4845 ( .IN1(\read_value_mux[25][6] ), .IN2(n1631), .IN3(
        write_data[6]), .IN4(n3166), .Q(\words[25]/data_i[6] ) );
  AO22X1 U4846 ( .IN1(\read_value_mux[25][7] ), .IN2(n1631), .IN3(
        write_data[7]), .IN4(n3166), .Q(\words[25]/data_i[7] ) );
  AO22X1 U4847 ( .IN1(\read_value_mux[25][8] ), .IN2(n1631), .IN3(
        write_data[8]), .IN4(n3166), .Q(\words[25]/data_i[8] ) );
  AO22X1 U4848 ( .IN1(\read_value_mux[25][9] ), .IN2(n1631), .IN3(
        write_data[9]), .IN4(n3166), .Q(\words[25]/data_i[9] ) );
  AO21X1 U4849 ( .IN1(\words[25]/valid_o ), .IN2(n1743), .IN3(n3166), .Q(
        \words[25]/valid_i ) );
  AO22X1 U4850 ( .IN1(\read_value_mux[26][0] ), .IN2(n1639), .IN3(
        write_data[0]), .IN4(n3167), .Q(\words[26]/data_i[0] ) );
  AO22X1 U4851 ( .IN1(\read_value_mux[26][10] ), .IN2(n1639), .IN3(
        write_data[10]), .IN4(n3167), .Q(\words[26]/data_i[10] ) );
  AO22X1 U4852 ( .IN1(\read_value_mux[26][11] ), .IN2(n1639), .IN3(
        write_data[11]), .IN4(n3167), .Q(\words[26]/data_i[11] ) );
  AO22X1 U4853 ( .IN1(\read_value_mux[26][12] ), .IN2(n1639), .IN3(
        write_data[12]), .IN4(n3167), .Q(\words[26]/data_i[12] ) );
  AO22X1 U4854 ( .IN1(\read_value_mux[26][13] ), .IN2(n1639), .IN3(
        write_data[13]), .IN4(n3167), .Q(\words[26]/data_i[13] ) );
  AO22X1 U4855 ( .IN1(\read_value_mux[26][14] ), .IN2(n1639), .IN3(
        write_data[14]), .IN4(n3167), .Q(\words[26]/data_i[14] ) );
  AO22X1 U4856 ( .IN1(\read_value_mux[26][15] ), .IN2(n1639), .IN3(
        write_data[15]), .IN4(n3167), .Q(\words[26]/data_i[15] ) );
  AO22X1 U4857 ( .IN1(\read_value_mux[26][16] ), .IN2(n1639), .IN3(
        write_data[16]), .IN4(n3167), .Q(\words[26]/data_i[16] ) );
  AO22X1 U4858 ( .IN1(\read_value_mux[26][17] ), .IN2(n1639), .IN3(
        write_data[17]), .IN4(n3167), .Q(\words[26]/data_i[17] ) );
  AO22X1 U4859 ( .IN1(\read_value_mux[26][18] ), .IN2(n1639), .IN3(
        write_data[18]), .IN4(n3167), .Q(\words[26]/data_i[18] ) );
  AO22X1 U4860 ( .IN1(\read_value_mux[26][19] ), .IN2(n1639), .IN3(
        write_data[19]), .IN4(n3167), .Q(\words[26]/data_i[19] ) );
  AO22X1 U4861 ( .IN1(\read_value_mux[26][1] ), .IN2(n1639), .IN3(
        write_data[1]), .IN4(n3167), .Q(\words[26]/data_i[1] ) );
  AO22X1 U4862 ( .IN1(\read_value_mux[26][20] ), .IN2(n1639), .IN3(
        write_data[20]), .IN4(n3167), .Q(\words[26]/data_i[20] ) );
  AO22X1 U4863 ( .IN1(\read_value_mux[26][21] ), .IN2(n1639), .IN3(
        write_data[21]), .IN4(n3167), .Q(\words[26]/data_i[21] ) );
  AO22X1 U4864 ( .IN1(\read_value_mux[26][22] ), .IN2(n1639), .IN3(
        write_data[22]), .IN4(n3167), .Q(\words[26]/data_i[22] ) );
  AO22X1 U4865 ( .IN1(\read_value_mux[26][23] ), .IN2(n1639), .IN3(
        write_data[23]), .IN4(n3167), .Q(\words[26]/data_i[23] ) );
  AO22X1 U4866 ( .IN1(\read_value_mux[26][24] ), .IN2(n1639), .IN3(
        write_data[24]), .IN4(n3167), .Q(\words[26]/data_i[24] ) );
  AO22X1 U4867 ( .IN1(\read_value_mux[26][25] ), .IN2(n1639), .IN3(
        write_data[25]), .IN4(n3167), .Q(\words[26]/data_i[25] ) );
  AO22X1 U4868 ( .IN1(\read_value_mux[26][26] ), .IN2(n1639), .IN3(
        write_data[26]), .IN4(n3167), .Q(\words[26]/data_i[26] ) );
  AO22X1 U4869 ( .IN1(\read_value_mux[26][27] ), .IN2(n1639), .IN3(
        write_data[27]), .IN4(n3167), .Q(\words[26]/data_i[27] ) );
  AO22X1 U4870 ( .IN1(\read_value_mux[26][28] ), .IN2(n1639), .IN3(
        write_data[28]), .IN4(n3167), .Q(\words[26]/data_i[28] ) );
  AO22X1 U4871 ( .IN1(\read_value_mux[26][29] ), .IN2(n1639), .IN3(
        write_data[29]), .IN4(n3167), .Q(\words[26]/data_i[29] ) );
  AO22X1 U4872 ( .IN1(\read_value_mux[26][2] ), .IN2(n1639), .IN3(
        write_data[2]), .IN4(n3167), .Q(\words[26]/data_i[2] ) );
  AO22X1 U4873 ( .IN1(\read_value_mux[26][30] ), .IN2(n1639), .IN3(
        write_data[30]), .IN4(n3167), .Q(\words[26]/data_i[30] ) );
  AO22X1 U4874 ( .IN1(\read_value_mux[26][31] ), .IN2(n1639), .IN3(
        write_data[31]), .IN4(n3167), .Q(\words[26]/data_i[31] ) );
  AO22X1 U4875 ( .IN1(\read_value_mux[26][3] ), .IN2(n1639), .IN3(
        write_data[3]), .IN4(n3167), .Q(\words[26]/data_i[3] ) );
  AO22X1 U4876 ( .IN1(\read_value_mux[26][4] ), .IN2(n1639), .IN3(
        write_data[4]), .IN4(n3167), .Q(\words[26]/data_i[4] ) );
  AO22X1 U4877 ( .IN1(\read_value_mux[26][5] ), .IN2(n1639), .IN3(
        write_data[5]), .IN4(n3167), .Q(\words[26]/data_i[5] ) );
  AO22X1 U4878 ( .IN1(\read_value_mux[26][6] ), .IN2(n1639), .IN3(
        write_data[6]), .IN4(n3167), .Q(\words[26]/data_i[6] ) );
  AO22X1 U4879 ( .IN1(\read_value_mux[26][7] ), .IN2(n1639), .IN3(
        write_data[7]), .IN4(n3167), .Q(\words[26]/data_i[7] ) );
  AO22X1 U4880 ( .IN1(\read_value_mux[26][8] ), .IN2(n1639), .IN3(
        write_data[8]), .IN4(n3167), .Q(\words[26]/data_i[8] ) );
  AO22X1 U4881 ( .IN1(\read_value_mux[26][9] ), .IN2(n1639), .IN3(
        write_data[9]), .IN4(n3167), .Q(\words[26]/data_i[9] ) );
  AO21X1 U4882 ( .IN1(\words[26]/valid_o ), .IN2(n1743), .IN3(n3167), .Q(
        \words[26]/valid_i ) );
  AO22X1 U4883 ( .IN1(\read_value_mux[27][0] ), .IN2(n1640), .IN3(
        write_data[0]), .IN4(n3169), .Q(\words[27]/data_i[0] ) );
  AO22X1 U4884 ( .IN1(\read_value_mux[27][10] ), .IN2(n1640), .IN3(
        write_data[10]), .IN4(n3169), .Q(\words[27]/data_i[10] ) );
  AO22X1 U4885 ( .IN1(\read_value_mux[27][11] ), .IN2(n1640), .IN3(
        write_data[11]), .IN4(n3169), .Q(\words[27]/data_i[11] ) );
  AO22X1 U4886 ( .IN1(\read_value_mux[27][12] ), .IN2(n1640), .IN3(
        write_data[12]), .IN4(n3169), .Q(\words[27]/data_i[12] ) );
  AO22X1 U4887 ( .IN1(\read_value_mux[27][13] ), .IN2(n1640), .IN3(
        write_data[13]), .IN4(n3169), .Q(\words[27]/data_i[13] ) );
  AO22X1 U4888 ( .IN1(\read_value_mux[27][14] ), .IN2(n1640), .IN3(
        write_data[14]), .IN4(n3169), .Q(\words[27]/data_i[14] ) );
  AO22X1 U4889 ( .IN1(\read_value_mux[27][15] ), .IN2(n1640), .IN3(
        write_data[15]), .IN4(n3169), .Q(\words[27]/data_i[15] ) );
  AO22X1 U4890 ( .IN1(\read_value_mux[27][16] ), .IN2(n1640), .IN3(
        write_data[16]), .IN4(n3169), .Q(\words[27]/data_i[16] ) );
  AO22X1 U4891 ( .IN1(\read_value_mux[27][17] ), .IN2(n1640), .IN3(
        write_data[17]), .IN4(n3169), .Q(\words[27]/data_i[17] ) );
  AO22X1 U4892 ( .IN1(\read_value_mux[27][18] ), .IN2(n1640), .IN3(
        write_data[18]), .IN4(n3169), .Q(\words[27]/data_i[18] ) );
  AO22X1 U4893 ( .IN1(\read_value_mux[27][19] ), .IN2(n1640), .IN3(
        write_data[19]), .IN4(n3169), .Q(\words[27]/data_i[19] ) );
  AO22X1 U4894 ( .IN1(\read_value_mux[27][1] ), .IN2(n1640), .IN3(
        write_data[1]), .IN4(n3169), .Q(\words[27]/data_i[1] ) );
  AO22X1 U4895 ( .IN1(\read_value_mux[27][20] ), .IN2(n1640), .IN3(
        write_data[20]), .IN4(n3169), .Q(\words[27]/data_i[20] ) );
  AO22X1 U4896 ( .IN1(\read_value_mux[27][21] ), .IN2(n1640), .IN3(
        write_data[21]), .IN4(n3169), .Q(\words[27]/data_i[21] ) );
  AO22X1 U4897 ( .IN1(\read_value_mux[27][22] ), .IN2(n1640), .IN3(
        write_data[22]), .IN4(n3169), .Q(\words[27]/data_i[22] ) );
  AO22X1 U4898 ( .IN1(\read_value_mux[27][23] ), .IN2(n1640), .IN3(
        write_data[23]), .IN4(n3169), .Q(\words[27]/data_i[23] ) );
  AO22X1 U4899 ( .IN1(\read_value_mux[27][24] ), .IN2(n1640), .IN3(
        write_data[24]), .IN4(n3169), .Q(\words[27]/data_i[24] ) );
  AO22X1 U4900 ( .IN1(\read_value_mux[27][25] ), .IN2(n1640), .IN3(
        write_data[25]), .IN4(n3169), .Q(\words[27]/data_i[25] ) );
  AO22X1 U4901 ( .IN1(\read_value_mux[27][26] ), .IN2(n1640), .IN3(
        write_data[26]), .IN4(n3169), .Q(\words[27]/data_i[26] ) );
  AO22X1 U4902 ( .IN1(\read_value_mux[27][27] ), .IN2(n1640), .IN3(
        write_data[27]), .IN4(n3169), .Q(\words[27]/data_i[27] ) );
  AO22X1 U4903 ( .IN1(\read_value_mux[27][28] ), .IN2(n1640), .IN3(
        write_data[28]), .IN4(n3169), .Q(\words[27]/data_i[28] ) );
  AO22X1 U4904 ( .IN1(\read_value_mux[27][29] ), .IN2(n1640), .IN3(
        write_data[29]), .IN4(n3169), .Q(\words[27]/data_i[29] ) );
  AO22X1 U4905 ( .IN1(\read_value_mux[27][2] ), .IN2(n1640), .IN3(
        write_data[2]), .IN4(n3169), .Q(\words[27]/data_i[2] ) );
  AO22X1 U4906 ( .IN1(\read_value_mux[27][30] ), .IN2(n1640), .IN3(
        write_data[30]), .IN4(n3169), .Q(\words[27]/data_i[30] ) );
  AO22X1 U4907 ( .IN1(\read_value_mux[27][31] ), .IN2(n1640), .IN3(
        write_data[31]), .IN4(n3169), .Q(\words[27]/data_i[31] ) );
  AO22X1 U4908 ( .IN1(\read_value_mux[27][3] ), .IN2(n1640), .IN3(
        write_data[3]), .IN4(n3169), .Q(\words[27]/data_i[3] ) );
  AO22X1 U4909 ( .IN1(\read_value_mux[27][4] ), .IN2(n1640), .IN3(
        write_data[4]), .IN4(n3169), .Q(\words[27]/data_i[4] ) );
  AO22X1 U4910 ( .IN1(\read_value_mux[27][5] ), .IN2(n1640), .IN3(
        write_data[5]), .IN4(n3169), .Q(\words[27]/data_i[5] ) );
  AO22X1 U4911 ( .IN1(\read_value_mux[27][6] ), .IN2(n1640), .IN3(
        write_data[6]), .IN4(n3169), .Q(\words[27]/data_i[6] ) );
  AO22X1 U4912 ( .IN1(\read_value_mux[27][7] ), .IN2(n1640), .IN3(
        write_data[7]), .IN4(n3169), .Q(\words[27]/data_i[7] ) );
  AO22X1 U4913 ( .IN1(\read_value_mux[27][8] ), .IN2(n1640), .IN3(
        write_data[8]), .IN4(n3169), .Q(\words[27]/data_i[8] ) );
  AO22X1 U4914 ( .IN1(\read_value_mux[27][9] ), .IN2(n1640), .IN3(
        write_data[9]), .IN4(n3169), .Q(\words[27]/data_i[9] ) );
  AO21X1 U4915 ( .IN1(\words[27]/valid_o ), .IN2(n1743), .IN3(n3169), .Q(
        \words[27]/valid_i ) );
  AO22X1 U4916 ( .IN1(\read_value_mux[28][0] ), .IN2(n1632), .IN3(
        write_data[0]), .IN4(n3171), .Q(\words[28]/data_i[0] ) );
  AO22X1 U4917 ( .IN1(\read_value_mux[28][10] ), .IN2(n1632), .IN3(
        write_data[10]), .IN4(n3171), .Q(\words[28]/data_i[10] ) );
  AO22X1 U4918 ( .IN1(\read_value_mux[28][11] ), .IN2(n1632), .IN3(
        write_data[11]), .IN4(n3171), .Q(\words[28]/data_i[11] ) );
  AO22X1 U4919 ( .IN1(\read_value_mux[28][12] ), .IN2(n1632), .IN3(
        write_data[12]), .IN4(n3171), .Q(\words[28]/data_i[12] ) );
  AO22X1 U4920 ( .IN1(\read_value_mux[28][13] ), .IN2(n1632), .IN3(
        write_data[13]), .IN4(n3171), .Q(\words[28]/data_i[13] ) );
  AO22X1 U4921 ( .IN1(\read_value_mux[28][14] ), .IN2(n1632), .IN3(
        write_data[14]), .IN4(n3171), .Q(\words[28]/data_i[14] ) );
  AO22X1 U4922 ( .IN1(\read_value_mux[28][15] ), .IN2(n1632), .IN3(
        write_data[15]), .IN4(n3171), .Q(\words[28]/data_i[15] ) );
  AO22X1 U4923 ( .IN1(\read_value_mux[28][16] ), .IN2(n1632), .IN3(
        write_data[16]), .IN4(n3171), .Q(\words[28]/data_i[16] ) );
  AO22X1 U4924 ( .IN1(\read_value_mux[28][17] ), .IN2(n1632), .IN3(
        write_data[17]), .IN4(n3171), .Q(\words[28]/data_i[17] ) );
  AO22X1 U4925 ( .IN1(\read_value_mux[28][18] ), .IN2(n1632), .IN3(
        write_data[18]), .IN4(n3171), .Q(\words[28]/data_i[18] ) );
  AO22X1 U4926 ( .IN1(\read_value_mux[28][19] ), .IN2(n1632), .IN3(
        write_data[19]), .IN4(n3171), .Q(\words[28]/data_i[19] ) );
  AO22X1 U4927 ( .IN1(\read_value_mux[28][1] ), .IN2(n1632), .IN3(
        write_data[1]), .IN4(n3171), .Q(\words[28]/data_i[1] ) );
  AO22X1 U4928 ( .IN1(\read_value_mux[28][20] ), .IN2(n1632), .IN3(
        write_data[20]), .IN4(n3171), .Q(\words[28]/data_i[20] ) );
  AO22X1 U4929 ( .IN1(\read_value_mux[28][21] ), .IN2(n1632), .IN3(
        write_data[21]), .IN4(n3171), .Q(\words[28]/data_i[21] ) );
  AO22X1 U4930 ( .IN1(\read_value_mux[28][22] ), .IN2(n1632), .IN3(
        write_data[22]), .IN4(n3171), .Q(\words[28]/data_i[22] ) );
  AO22X1 U4931 ( .IN1(\read_value_mux[28][23] ), .IN2(n1632), .IN3(
        write_data[23]), .IN4(n3171), .Q(\words[28]/data_i[23] ) );
  AO22X1 U4932 ( .IN1(\read_value_mux[28][24] ), .IN2(n1632), .IN3(
        write_data[24]), .IN4(n3171), .Q(\words[28]/data_i[24] ) );
  AO22X1 U4933 ( .IN1(\read_value_mux[28][25] ), .IN2(n1632), .IN3(
        write_data[25]), .IN4(n3171), .Q(\words[28]/data_i[25] ) );
  AO22X1 U4934 ( .IN1(\read_value_mux[28][26] ), .IN2(n1632), .IN3(
        write_data[26]), .IN4(n3171), .Q(\words[28]/data_i[26] ) );
  AO22X1 U4935 ( .IN1(\read_value_mux[28][27] ), .IN2(n1632), .IN3(
        write_data[27]), .IN4(n3171), .Q(\words[28]/data_i[27] ) );
  AO22X1 U4936 ( .IN1(\read_value_mux[28][28] ), .IN2(n1632), .IN3(
        write_data[28]), .IN4(n3171), .Q(\words[28]/data_i[28] ) );
  AO22X1 U4937 ( .IN1(\read_value_mux[28][29] ), .IN2(n1632), .IN3(
        write_data[29]), .IN4(n3171), .Q(\words[28]/data_i[29] ) );
  AO22X1 U4938 ( .IN1(\read_value_mux[28][2] ), .IN2(n1632), .IN3(
        write_data[2]), .IN4(n3171), .Q(\words[28]/data_i[2] ) );
  AO22X1 U4939 ( .IN1(\read_value_mux[28][30] ), .IN2(n1632), .IN3(
        write_data[30]), .IN4(n3171), .Q(\words[28]/data_i[30] ) );
  AO22X1 U4940 ( .IN1(\read_value_mux[28][31] ), .IN2(n1632), .IN3(
        write_data[31]), .IN4(n3171), .Q(\words[28]/data_i[31] ) );
  AO22X1 U4941 ( .IN1(\read_value_mux[28][3] ), .IN2(n1632), .IN3(
        write_data[3]), .IN4(n3171), .Q(\words[28]/data_i[3] ) );
  AO22X1 U4942 ( .IN1(\read_value_mux[28][4] ), .IN2(n1632), .IN3(
        write_data[4]), .IN4(n3171), .Q(\words[28]/data_i[4] ) );
  AO22X1 U4943 ( .IN1(\read_value_mux[28][5] ), .IN2(n1632), .IN3(
        write_data[5]), .IN4(n3171), .Q(\words[28]/data_i[5] ) );
  AO22X1 U4944 ( .IN1(\read_value_mux[28][6] ), .IN2(n1632), .IN3(
        write_data[6]), .IN4(n3171), .Q(\words[28]/data_i[6] ) );
  AO22X1 U4945 ( .IN1(\read_value_mux[28][7] ), .IN2(n1632), .IN3(
        write_data[7]), .IN4(n3171), .Q(\words[28]/data_i[7] ) );
  AO22X1 U4946 ( .IN1(\read_value_mux[28][8] ), .IN2(n1632), .IN3(
        write_data[8]), .IN4(n3171), .Q(\words[28]/data_i[8] ) );
  AO22X1 U4947 ( .IN1(\read_value_mux[28][9] ), .IN2(n1632), .IN3(
        write_data[9]), .IN4(n3171), .Q(\words[28]/data_i[9] ) );
  AO21X1 U4948 ( .IN1(\words[28]/valid_o ), .IN2(n1743), .IN3(n3171), .Q(
        \words[28]/valid_i ) );
  AO22X1 U4949 ( .IN1(\read_value_mux[29][0] ), .IN2(n1633), .IN3(
        write_data[0]), .IN4(n3172), .Q(\words[29]/data_i[0] ) );
  AO22X1 U4950 ( .IN1(\read_value_mux[29][10] ), .IN2(n1633), .IN3(
        write_data[10]), .IN4(n3172), .Q(\words[29]/data_i[10] ) );
  AO22X1 U4951 ( .IN1(\read_value_mux[29][11] ), .IN2(n1633), .IN3(
        write_data[11]), .IN4(n3172), .Q(\words[29]/data_i[11] ) );
  AO22X1 U4952 ( .IN1(\read_value_mux[29][12] ), .IN2(n1633), .IN3(
        write_data[12]), .IN4(n3172), .Q(\words[29]/data_i[12] ) );
  AO22X1 U4953 ( .IN1(\read_value_mux[29][13] ), .IN2(n1633), .IN3(
        write_data[13]), .IN4(n3172), .Q(\words[29]/data_i[13] ) );
  AO22X1 U4954 ( .IN1(\read_value_mux[29][14] ), .IN2(n1633), .IN3(
        write_data[14]), .IN4(n3172), .Q(\words[29]/data_i[14] ) );
  AO22X1 U4955 ( .IN1(\read_value_mux[29][15] ), .IN2(n1633), .IN3(
        write_data[15]), .IN4(n3172), .Q(\words[29]/data_i[15] ) );
  AO22X1 U4956 ( .IN1(\read_value_mux[29][16] ), .IN2(n1633), .IN3(
        write_data[16]), .IN4(n3172), .Q(\words[29]/data_i[16] ) );
  AO22X1 U4957 ( .IN1(\read_value_mux[29][17] ), .IN2(n1633), .IN3(
        write_data[17]), .IN4(n3172), .Q(\words[29]/data_i[17] ) );
  AO22X1 U4958 ( .IN1(\read_value_mux[29][18] ), .IN2(n1633), .IN3(
        write_data[18]), .IN4(n3172), .Q(\words[29]/data_i[18] ) );
  AO22X1 U4959 ( .IN1(\read_value_mux[29][19] ), .IN2(n1633), .IN3(
        write_data[19]), .IN4(n3172), .Q(\words[29]/data_i[19] ) );
  AO22X1 U4960 ( .IN1(\read_value_mux[29][1] ), .IN2(n1633), .IN3(
        write_data[1]), .IN4(n3172), .Q(\words[29]/data_i[1] ) );
  AO22X1 U4961 ( .IN1(\read_value_mux[29][20] ), .IN2(n1633), .IN3(
        write_data[20]), .IN4(n3172), .Q(\words[29]/data_i[20] ) );
  AO22X1 U4962 ( .IN1(\read_value_mux[29][21] ), .IN2(n1633), .IN3(
        write_data[21]), .IN4(n3172), .Q(\words[29]/data_i[21] ) );
  AO22X1 U4963 ( .IN1(\read_value_mux[29][22] ), .IN2(n1633), .IN3(
        write_data[22]), .IN4(n3172), .Q(\words[29]/data_i[22] ) );
  AO22X1 U4964 ( .IN1(\read_value_mux[29][23] ), .IN2(n1633), .IN3(
        write_data[23]), .IN4(n3172), .Q(\words[29]/data_i[23] ) );
  AO22X1 U4965 ( .IN1(\read_value_mux[29][24] ), .IN2(n1633), .IN3(
        write_data[24]), .IN4(n3172), .Q(\words[29]/data_i[24] ) );
  AO22X1 U4966 ( .IN1(\read_value_mux[29][25] ), .IN2(n1633), .IN3(
        write_data[25]), .IN4(n3172), .Q(\words[29]/data_i[25] ) );
  AO22X1 U4967 ( .IN1(\read_value_mux[29][26] ), .IN2(n1633), .IN3(
        write_data[26]), .IN4(n3172), .Q(\words[29]/data_i[26] ) );
  AO22X1 U4968 ( .IN1(\read_value_mux[29][27] ), .IN2(n1633), .IN3(
        write_data[27]), .IN4(n3172), .Q(\words[29]/data_i[27] ) );
  AO22X1 U4969 ( .IN1(\read_value_mux[29][28] ), .IN2(n1633), .IN3(
        write_data[28]), .IN4(n3172), .Q(\words[29]/data_i[28] ) );
  AO22X1 U4970 ( .IN1(\read_value_mux[29][29] ), .IN2(n1633), .IN3(
        write_data[29]), .IN4(n3172), .Q(\words[29]/data_i[29] ) );
  AO22X1 U4971 ( .IN1(\read_value_mux[29][2] ), .IN2(n1633), .IN3(
        write_data[2]), .IN4(n3172), .Q(\words[29]/data_i[2] ) );
  AO22X1 U4972 ( .IN1(\read_value_mux[29][30] ), .IN2(n1633), .IN3(
        write_data[30]), .IN4(n3172), .Q(\words[29]/data_i[30] ) );
  AO22X1 U4973 ( .IN1(\read_value_mux[29][31] ), .IN2(n1633), .IN3(
        write_data[31]), .IN4(n3172), .Q(\words[29]/data_i[31] ) );
  AO22X1 U4974 ( .IN1(\read_value_mux[29][3] ), .IN2(n1633), .IN3(
        write_data[3]), .IN4(n3172), .Q(\words[29]/data_i[3] ) );
  AO22X1 U4975 ( .IN1(\read_value_mux[29][4] ), .IN2(n1633), .IN3(
        write_data[4]), .IN4(n3172), .Q(\words[29]/data_i[4] ) );
  AO22X1 U4976 ( .IN1(\read_value_mux[29][5] ), .IN2(n1633), .IN3(
        write_data[5]), .IN4(n3172), .Q(\words[29]/data_i[5] ) );
  AO22X1 U4977 ( .IN1(\read_value_mux[29][6] ), .IN2(n1633), .IN3(
        write_data[6]), .IN4(n3172), .Q(\words[29]/data_i[6] ) );
  AO22X1 U4978 ( .IN1(\read_value_mux[29][7] ), .IN2(n1633), .IN3(
        write_data[7]), .IN4(n3172), .Q(\words[29]/data_i[7] ) );
  AO22X1 U4979 ( .IN1(\read_value_mux[29][8] ), .IN2(n1633), .IN3(
        write_data[8]), .IN4(n3172), .Q(\words[29]/data_i[8] ) );
  AO22X1 U4980 ( .IN1(\read_value_mux[29][9] ), .IN2(n1633), .IN3(
        write_data[9]), .IN4(n3172), .Q(\words[29]/data_i[9] ) );
  AO21X1 U4981 ( .IN1(\words[29]/valid_o ), .IN2(n1743), .IN3(n3172), .Q(
        \words[29]/valid_i ) );
  AO22X1 U4982 ( .IN1(\read_value_mux[2][0] ), .IN2(n1615), .IN3(write_data[0]), .IN4(n3173), .Q(\words[2]/data_i[0] ) );
  AO22X1 U4983 ( .IN1(\read_value_mux[2][10] ), .IN2(n1615), .IN3(
        write_data[10]), .IN4(n3173), .Q(\words[2]/data_i[10] ) );
  AO22X1 U4984 ( .IN1(\read_value_mux[2][11] ), .IN2(n1615), .IN3(
        write_data[11]), .IN4(n3173), .Q(\words[2]/data_i[11] ) );
  AO22X1 U4985 ( .IN1(\read_value_mux[2][12] ), .IN2(n1615), .IN3(
        write_data[12]), .IN4(n3173), .Q(\words[2]/data_i[12] ) );
  AO22X1 U4986 ( .IN1(\read_value_mux[2][13] ), .IN2(n1615), .IN3(
        write_data[13]), .IN4(n3173), .Q(\words[2]/data_i[13] ) );
  AO22X1 U4987 ( .IN1(\read_value_mux[2][14] ), .IN2(n1615), .IN3(
        write_data[14]), .IN4(n3173), .Q(\words[2]/data_i[14] ) );
  AO22X1 U4988 ( .IN1(\read_value_mux[2][15] ), .IN2(n1615), .IN3(
        write_data[15]), .IN4(n3173), .Q(\words[2]/data_i[15] ) );
  AO22X1 U4989 ( .IN1(\read_value_mux[2][16] ), .IN2(n1615), .IN3(
        write_data[16]), .IN4(n3173), .Q(\words[2]/data_i[16] ) );
  AO22X1 U4990 ( .IN1(\read_value_mux[2][17] ), .IN2(n1615), .IN3(
        write_data[17]), .IN4(n3173), .Q(\words[2]/data_i[17] ) );
  AO22X1 U4991 ( .IN1(\read_value_mux[2][18] ), .IN2(n1615), .IN3(
        write_data[18]), .IN4(n3173), .Q(\words[2]/data_i[18] ) );
  AO22X1 U4992 ( .IN1(\read_value_mux[2][19] ), .IN2(n1615), .IN3(
        write_data[19]), .IN4(n3173), .Q(\words[2]/data_i[19] ) );
  AO22X1 U4993 ( .IN1(\read_value_mux[2][1] ), .IN2(n1615), .IN3(write_data[1]), .IN4(n3173), .Q(\words[2]/data_i[1] ) );
  AO22X1 U4994 ( .IN1(\read_value_mux[2][20] ), .IN2(n1615), .IN3(
        write_data[20]), .IN4(n3173), .Q(\words[2]/data_i[20] ) );
  AO22X1 U4995 ( .IN1(\read_value_mux[2][21] ), .IN2(n1615), .IN3(
        write_data[21]), .IN4(n3173), .Q(\words[2]/data_i[21] ) );
  AO22X1 U4996 ( .IN1(\read_value_mux[2][22] ), .IN2(n1615), .IN3(
        write_data[22]), .IN4(n3173), .Q(\words[2]/data_i[22] ) );
  AO22X1 U4997 ( .IN1(\read_value_mux[2][23] ), .IN2(n1615), .IN3(
        write_data[23]), .IN4(n3173), .Q(\words[2]/data_i[23] ) );
  AO22X1 U4998 ( .IN1(\read_value_mux[2][24] ), .IN2(n1615), .IN3(
        write_data[24]), .IN4(n3173), .Q(\words[2]/data_i[24] ) );
  AO22X1 U4999 ( .IN1(\read_value_mux[2][25] ), .IN2(n1615), .IN3(
        write_data[25]), .IN4(n3173), .Q(\words[2]/data_i[25] ) );
  AO22X1 U5000 ( .IN1(\read_value_mux[2][26] ), .IN2(n1615), .IN3(
        write_data[26]), .IN4(n3173), .Q(\words[2]/data_i[26] ) );
  AO22X1 U5001 ( .IN1(\read_value_mux[2][27] ), .IN2(n1615), .IN3(
        write_data[27]), .IN4(n3173), .Q(\words[2]/data_i[27] ) );
  AO22X1 U5002 ( .IN1(\read_value_mux[2][28] ), .IN2(n1615), .IN3(
        write_data[28]), .IN4(n3173), .Q(\words[2]/data_i[28] ) );
  AO22X1 U5003 ( .IN1(\read_value_mux[2][29] ), .IN2(n1615), .IN3(
        write_data[29]), .IN4(n3173), .Q(\words[2]/data_i[29] ) );
  AO22X1 U5004 ( .IN1(\read_value_mux[2][2] ), .IN2(n1615), .IN3(write_data[2]), .IN4(n3173), .Q(\words[2]/data_i[2] ) );
  AO22X1 U5005 ( .IN1(\read_value_mux[2][30] ), .IN2(n1615), .IN3(
        write_data[30]), .IN4(n3173), .Q(\words[2]/data_i[30] ) );
  AO22X1 U5006 ( .IN1(\read_value_mux[2][31] ), .IN2(n1615), .IN3(
        write_data[31]), .IN4(n3173), .Q(\words[2]/data_i[31] ) );
  AO22X1 U5007 ( .IN1(\read_value_mux[2][3] ), .IN2(n1615), .IN3(write_data[3]), .IN4(n3173), .Q(\words[2]/data_i[3] ) );
  AO22X1 U5008 ( .IN1(\read_value_mux[2][4] ), .IN2(n1615), .IN3(write_data[4]), .IN4(n3173), .Q(\words[2]/data_i[4] ) );
  AO22X1 U5009 ( .IN1(\read_value_mux[2][5] ), .IN2(n1615), .IN3(write_data[5]), .IN4(n3173), .Q(\words[2]/data_i[5] ) );
  AO22X1 U5010 ( .IN1(\read_value_mux[2][6] ), .IN2(n1615), .IN3(write_data[6]), .IN4(n3173), .Q(\words[2]/data_i[6] ) );
  AO22X1 U5011 ( .IN1(\read_value_mux[2][7] ), .IN2(n1615), .IN3(write_data[7]), .IN4(n3173), .Q(\words[2]/data_i[7] ) );
  AO22X1 U5012 ( .IN1(\read_value_mux[2][8] ), .IN2(n1615), .IN3(write_data[8]), .IN4(n3173), .Q(\words[2]/data_i[8] ) );
  AO22X1 U5013 ( .IN1(\read_value_mux[2][9] ), .IN2(n1615), .IN3(write_data[9]), .IN4(n3173), .Q(\words[2]/data_i[9] ) );
  AO21X1 U5014 ( .IN1(\words[2]/valid_o ), .IN2(n1743), .IN3(n3173), .Q(
        \words[2]/valid_i ) );
  AO22X1 U5015 ( .IN1(\read_value_mux[30][0] ), .IN2(n1641), .IN3(
        write_data[0]), .IN4(n3174), .Q(\words[30]/data_i[0] ) );
  AO22X1 U5016 ( .IN1(\read_value_mux[30][10] ), .IN2(n1641), .IN3(
        write_data[10]), .IN4(n3174), .Q(\words[30]/data_i[10] ) );
  AO22X1 U5017 ( .IN1(\read_value_mux[30][11] ), .IN2(n1641), .IN3(
        write_data[11]), .IN4(n3174), .Q(\words[30]/data_i[11] ) );
  AO22X1 U5018 ( .IN1(\read_value_mux[30][12] ), .IN2(n1641), .IN3(
        write_data[12]), .IN4(n3174), .Q(\words[30]/data_i[12] ) );
  AO22X1 U5019 ( .IN1(\read_value_mux[30][13] ), .IN2(n1641), .IN3(
        write_data[13]), .IN4(n3174), .Q(\words[30]/data_i[13] ) );
  AO22X1 U5020 ( .IN1(\read_value_mux[30][14] ), .IN2(n1641), .IN3(
        write_data[14]), .IN4(n3174), .Q(\words[30]/data_i[14] ) );
  AO22X1 U5021 ( .IN1(\read_value_mux[30][15] ), .IN2(n1641), .IN3(
        write_data[15]), .IN4(n3174), .Q(\words[30]/data_i[15] ) );
  AO22X1 U5022 ( .IN1(\read_value_mux[30][16] ), .IN2(n1641), .IN3(
        write_data[16]), .IN4(n3174), .Q(\words[30]/data_i[16] ) );
  AO22X1 U5023 ( .IN1(\read_value_mux[30][17] ), .IN2(n1641), .IN3(
        write_data[17]), .IN4(n3174), .Q(\words[30]/data_i[17] ) );
  AO22X1 U5024 ( .IN1(\read_value_mux[30][18] ), .IN2(n1641), .IN3(
        write_data[18]), .IN4(n3174), .Q(\words[30]/data_i[18] ) );
  AO22X1 U5025 ( .IN1(\read_value_mux[30][19] ), .IN2(n1641), .IN3(
        write_data[19]), .IN4(n3174), .Q(\words[30]/data_i[19] ) );
  AO22X1 U5026 ( .IN1(\read_value_mux[30][1] ), .IN2(n1641), .IN3(
        write_data[1]), .IN4(n3174), .Q(\words[30]/data_i[1] ) );
  AO22X1 U5027 ( .IN1(\read_value_mux[30][20] ), .IN2(n1641), .IN3(
        write_data[20]), .IN4(n3174), .Q(\words[30]/data_i[20] ) );
  AO22X1 U5028 ( .IN1(\read_value_mux[30][21] ), .IN2(n1641), .IN3(
        write_data[21]), .IN4(n3174), .Q(\words[30]/data_i[21] ) );
  AO22X1 U5029 ( .IN1(\read_value_mux[30][22] ), .IN2(n1641), .IN3(
        write_data[22]), .IN4(n3174), .Q(\words[30]/data_i[22] ) );
  AO22X1 U5030 ( .IN1(\read_value_mux[30][23] ), .IN2(n1641), .IN3(
        write_data[23]), .IN4(n3174), .Q(\words[30]/data_i[23] ) );
  AO22X1 U5031 ( .IN1(\read_value_mux[30][24] ), .IN2(n1641), .IN3(
        write_data[24]), .IN4(n3174), .Q(\words[30]/data_i[24] ) );
  AO22X1 U5032 ( .IN1(\read_value_mux[30][25] ), .IN2(n1641), .IN3(
        write_data[25]), .IN4(n3174), .Q(\words[30]/data_i[25] ) );
  AO22X1 U5033 ( .IN1(\read_value_mux[30][26] ), .IN2(n1641), .IN3(
        write_data[26]), .IN4(n3174), .Q(\words[30]/data_i[26] ) );
  AO22X1 U5034 ( .IN1(\read_value_mux[30][27] ), .IN2(n1641), .IN3(
        write_data[27]), .IN4(n3174), .Q(\words[30]/data_i[27] ) );
  AO22X1 U5035 ( .IN1(\read_value_mux[30][28] ), .IN2(n1641), .IN3(
        write_data[28]), .IN4(n3174), .Q(\words[30]/data_i[28] ) );
  AO22X1 U5036 ( .IN1(\read_value_mux[30][29] ), .IN2(n1641), .IN3(
        write_data[29]), .IN4(n3174), .Q(\words[30]/data_i[29] ) );
  AO22X1 U5037 ( .IN1(\read_value_mux[30][2] ), .IN2(n1641), .IN3(
        write_data[2]), .IN4(n3174), .Q(\words[30]/data_i[2] ) );
  AO22X1 U5038 ( .IN1(\read_value_mux[30][30] ), .IN2(n1641), .IN3(
        write_data[30]), .IN4(n3174), .Q(\words[30]/data_i[30] ) );
  AO22X1 U5039 ( .IN1(\read_value_mux[30][31] ), .IN2(n1641), .IN3(
        write_data[31]), .IN4(n3174), .Q(\words[30]/data_i[31] ) );
  AO22X1 U5040 ( .IN1(\read_value_mux[30][3] ), .IN2(n1641), .IN3(
        write_data[3]), .IN4(n3174), .Q(\words[30]/data_i[3] ) );
  AO22X1 U5041 ( .IN1(\read_value_mux[30][4] ), .IN2(n1641), .IN3(
        write_data[4]), .IN4(n3174), .Q(\words[30]/data_i[4] ) );
  AO22X1 U5042 ( .IN1(\read_value_mux[30][5] ), .IN2(n1641), .IN3(
        write_data[5]), .IN4(n3174), .Q(\words[30]/data_i[5] ) );
  AO22X1 U5043 ( .IN1(\read_value_mux[30][6] ), .IN2(n1641), .IN3(
        write_data[6]), .IN4(n3174), .Q(\words[30]/data_i[6] ) );
  AO22X1 U5044 ( .IN1(\read_value_mux[30][7] ), .IN2(n1641), .IN3(
        write_data[7]), .IN4(n3174), .Q(\words[30]/data_i[7] ) );
  AO22X1 U5045 ( .IN1(\read_value_mux[30][8] ), .IN2(n1641), .IN3(
        write_data[8]), .IN4(n3174), .Q(\words[30]/data_i[8] ) );
  AO22X1 U5046 ( .IN1(\read_value_mux[30][9] ), .IN2(n1641), .IN3(
        write_data[9]), .IN4(n3174), .Q(\words[30]/data_i[9] ) );
  AO21X1 U5047 ( .IN1(\words[30]/valid_o ), .IN2(n1743), .IN3(n3174), .Q(
        \words[30]/valid_i ) );
  AO22X1 U5048 ( .IN1(\read_value_mux[31][0] ), .IN2(n1642), .IN3(
        write_data[0]), .IN4(n3176), .Q(\words[31]/data_i[0] ) );
  AO22X1 U5049 ( .IN1(\read_value_mux[31][10] ), .IN2(n1642), .IN3(
        write_data[10]), .IN4(n3176), .Q(\words[31]/data_i[10] ) );
  AO22X1 U5050 ( .IN1(\read_value_mux[31][11] ), .IN2(n1642), .IN3(
        write_data[11]), .IN4(n3176), .Q(\words[31]/data_i[11] ) );
  AO22X1 U5051 ( .IN1(\read_value_mux[31][12] ), .IN2(n1642), .IN3(
        write_data[12]), .IN4(n3176), .Q(\words[31]/data_i[12] ) );
  AO22X1 U5052 ( .IN1(\read_value_mux[31][13] ), .IN2(n1642), .IN3(
        write_data[13]), .IN4(n3176), .Q(\words[31]/data_i[13] ) );
  AO22X1 U5053 ( .IN1(\read_value_mux[31][14] ), .IN2(n1642), .IN3(
        write_data[14]), .IN4(n3176), .Q(\words[31]/data_i[14] ) );
  AO22X1 U5054 ( .IN1(\read_value_mux[31][15] ), .IN2(n1642), .IN3(
        write_data[15]), .IN4(n3176), .Q(\words[31]/data_i[15] ) );
  AO22X1 U5055 ( .IN1(\read_value_mux[31][16] ), .IN2(n1642), .IN3(
        write_data[16]), .IN4(n3176), .Q(\words[31]/data_i[16] ) );
  AO22X1 U5056 ( .IN1(\read_value_mux[31][17] ), .IN2(n1642), .IN3(
        write_data[17]), .IN4(n3176), .Q(\words[31]/data_i[17] ) );
  AO22X1 U5057 ( .IN1(\read_value_mux[31][18] ), .IN2(n1642), .IN3(
        write_data[18]), .IN4(n3176), .Q(\words[31]/data_i[18] ) );
  AO22X1 U5058 ( .IN1(\read_value_mux[31][19] ), .IN2(n1642), .IN3(
        write_data[19]), .IN4(n3176), .Q(\words[31]/data_i[19] ) );
  AO22X1 U5059 ( .IN1(\read_value_mux[31][1] ), .IN2(n1642), .IN3(
        write_data[1]), .IN4(n3176), .Q(\words[31]/data_i[1] ) );
  AO22X1 U5060 ( .IN1(\read_value_mux[31][20] ), .IN2(n1642), .IN3(
        write_data[20]), .IN4(n3176), .Q(\words[31]/data_i[20] ) );
  AO22X1 U5061 ( .IN1(\read_value_mux[31][21] ), .IN2(n1642), .IN3(
        write_data[21]), .IN4(n3176), .Q(\words[31]/data_i[21] ) );
  AO22X1 U5062 ( .IN1(\read_value_mux[31][22] ), .IN2(n1642), .IN3(
        write_data[22]), .IN4(n3176), .Q(\words[31]/data_i[22] ) );
  AO22X1 U5063 ( .IN1(\read_value_mux[31][23] ), .IN2(n1642), .IN3(
        write_data[23]), .IN4(n3176), .Q(\words[31]/data_i[23] ) );
  AO22X1 U5064 ( .IN1(\read_value_mux[31][24] ), .IN2(n1642), .IN3(
        write_data[24]), .IN4(n3176), .Q(\words[31]/data_i[24] ) );
  AO22X1 U5065 ( .IN1(\read_value_mux[31][25] ), .IN2(n1642), .IN3(
        write_data[25]), .IN4(n3176), .Q(\words[31]/data_i[25] ) );
  AO22X1 U5066 ( .IN1(\read_value_mux[31][26] ), .IN2(n1642), .IN3(
        write_data[26]), .IN4(n3176), .Q(\words[31]/data_i[26] ) );
  AO22X1 U5067 ( .IN1(\read_value_mux[31][27] ), .IN2(n1642), .IN3(
        write_data[27]), .IN4(n3176), .Q(\words[31]/data_i[27] ) );
  AO22X1 U5068 ( .IN1(\read_value_mux[31][28] ), .IN2(n1642), .IN3(
        write_data[28]), .IN4(n3176), .Q(\words[31]/data_i[28] ) );
  AO22X1 U5069 ( .IN1(\read_value_mux[31][29] ), .IN2(n1642), .IN3(
        write_data[29]), .IN4(n3176), .Q(\words[31]/data_i[29] ) );
  AO22X1 U5070 ( .IN1(\read_value_mux[31][2] ), .IN2(n1642), .IN3(
        write_data[2]), .IN4(n3176), .Q(\words[31]/data_i[2] ) );
  AO22X1 U5071 ( .IN1(\read_value_mux[31][30] ), .IN2(n1642), .IN3(
        write_data[30]), .IN4(n3176), .Q(\words[31]/data_i[30] ) );
  AO22X1 U5072 ( .IN1(\read_value_mux[31][31] ), .IN2(n1642), .IN3(
        write_data[31]), .IN4(n3176), .Q(\words[31]/data_i[31] ) );
  AO22X1 U5073 ( .IN1(\read_value_mux[31][3] ), .IN2(n1642), .IN3(
        write_data[3]), .IN4(n3176), .Q(\words[31]/data_i[3] ) );
  AO22X1 U5074 ( .IN1(\read_value_mux[31][4] ), .IN2(n1642), .IN3(
        write_data[4]), .IN4(n3176), .Q(\words[31]/data_i[4] ) );
  AO22X1 U5075 ( .IN1(\read_value_mux[31][5] ), .IN2(n1642), .IN3(
        write_data[5]), .IN4(n3176), .Q(\words[31]/data_i[5] ) );
  AO22X1 U5076 ( .IN1(\read_value_mux[31][6] ), .IN2(n1642), .IN3(
        write_data[6]), .IN4(n3176), .Q(\words[31]/data_i[6] ) );
  AO22X1 U5077 ( .IN1(\read_value_mux[31][7] ), .IN2(n1642), .IN3(
        write_data[7]), .IN4(n3176), .Q(\words[31]/data_i[7] ) );
  AO22X1 U5078 ( .IN1(\read_value_mux[31][8] ), .IN2(n1642), .IN3(
        write_data[8]), .IN4(n3176), .Q(\words[31]/data_i[8] ) );
  AO22X1 U5079 ( .IN1(\read_value_mux[31][9] ), .IN2(n1642), .IN3(
        write_data[9]), .IN4(n3176), .Q(\words[31]/data_i[9] ) );
  AO21X1 U5080 ( .IN1(\words[31]/valid_o ), .IN2(n1743), .IN3(n3176), .Q(
        \words[31]/valid_i ) );
  AO22X1 U5081 ( .IN1(\read_value_mux[3][0] ), .IN2(n1643), .IN3(write_data[0]), .IN4(n3178), .Q(\words[3]/data_i[0] ) );
  AO22X1 U5082 ( .IN1(\read_value_mux[3][10] ), .IN2(n1643), .IN3(
        write_data[10]), .IN4(n3178), .Q(\words[3]/data_i[10] ) );
  AO22X1 U5083 ( .IN1(\read_value_mux[3][11] ), .IN2(n1643), .IN3(
        write_data[11]), .IN4(n3178), .Q(\words[3]/data_i[11] ) );
  AO22X1 U5084 ( .IN1(\read_value_mux[3][12] ), .IN2(n1643), .IN3(
        write_data[12]), .IN4(n3178), .Q(\words[3]/data_i[12] ) );
  AO22X1 U5085 ( .IN1(\read_value_mux[3][13] ), .IN2(n1643), .IN3(
        write_data[13]), .IN4(n3178), .Q(\words[3]/data_i[13] ) );
  AO22X1 U5086 ( .IN1(\read_value_mux[3][14] ), .IN2(n1643), .IN3(
        write_data[14]), .IN4(n3178), .Q(\words[3]/data_i[14] ) );
  AO22X1 U5087 ( .IN1(\read_value_mux[3][15] ), .IN2(n1643), .IN3(
        write_data[15]), .IN4(n3178), .Q(\words[3]/data_i[15] ) );
  AO22X1 U5088 ( .IN1(\read_value_mux[3][16] ), .IN2(n1643), .IN3(
        write_data[16]), .IN4(n3178), .Q(\words[3]/data_i[16] ) );
  AO22X1 U5089 ( .IN1(\read_value_mux[3][17] ), .IN2(n1643), .IN3(
        write_data[17]), .IN4(n3178), .Q(\words[3]/data_i[17] ) );
  AO22X1 U5090 ( .IN1(\read_value_mux[3][18] ), .IN2(n1643), .IN3(
        write_data[18]), .IN4(n3178), .Q(\words[3]/data_i[18] ) );
  AO22X1 U5091 ( .IN1(\read_value_mux[3][19] ), .IN2(n1643), .IN3(
        write_data[19]), .IN4(n3178), .Q(\words[3]/data_i[19] ) );
  AO22X1 U5092 ( .IN1(\read_value_mux[3][1] ), .IN2(n1643), .IN3(write_data[1]), .IN4(n3178), .Q(\words[3]/data_i[1] ) );
  AO22X1 U5093 ( .IN1(\read_value_mux[3][20] ), .IN2(n1643), .IN3(
        write_data[20]), .IN4(n3178), .Q(\words[3]/data_i[20] ) );
  AO22X1 U5094 ( .IN1(\read_value_mux[3][21] ), .IN2(n1643), .IN3(
        write_data[21]), .IN4(n3178), .Q(\words[3]/data_i[21] ) );
  AO22X1 U5095 ( .IN1(\read_value_mux[3][22] ), .IN2(n1643), .IN3(
        write_data[22]), .IN4(n3178), .Q(\words[3]/data_i[22] ) );
  AO22X1 U5096 ( .IN1(\read_value_mux[3][23] ), .IN2(n1643), .IN3(
        write_data[23]), .IN4(n3178), .Q(\words[3]/data_i[23] ) );
  AO22X1 U5097 ( .IN1(\read_value_mux[3][24] ), .IN2(n1643), .IN3(
        write_data[24]), .IN4(n3178), .Q(\words[3]/data_i[24] ) );
  AO22X1 U5098 ( .IN1(\read_value_mux[3][25] ), .IN2(n1643), .IN3(
        write_data[25]), .IN4(n3178), .Q(\words[3]/data_i[25] ) );
  AO22X1 U5099 ( .IN1(\read_value_mux[3][26] ), .IN2(n1643), .IN3(
        write_data[26]), .IN4(n3178), .Q(\words[3]/data_i[26] ) );
  AO22X1 U5100 ( .IN1(\read_value_mux[3][27] ), .IN2(n1643), .IN3(
        write_data[27]), .IN4(n3178), .Q(\words[3]/data_i[27] ) );
  AO22X1 U5101 ( .IN1(\read_value_mux[3][28] ), .IN2(n1643), .IN3(
        write_data[28]), .IN4(n3178), .Q(\words[3]/data_i[28] ) );
  AO22X1 U5102 ( .IN1(\read_value_mux[3][29] ), .IN2(n1643), .IN3(
        write_data[29]), .IN4(n3178), .Q(\words[3]/data_i[29] ) );
  AO22X1 U5103 ( .IN1(\read_value_mux[3][2] ), .IN2(n1643), .IN3(write_data[2]), .IN4(n3178), .Q(\words[3]/data_i[2] ) );
  AO22X1 U5104 ( .IN1(\read_value_mux[3][30] ), .IN2(n1643), .IN3(
        write_data[30]), .IN4(n3178), .Q(\words[3]/data_i[30] ) );
  AO22X1 U5105 ( .IN1(\read_value_mux[3][31] ), .IN2(n1643), .IN3(
        write_data[31]), .IN4(n3178), .Q(\words[3]/data_i[31] ) );
  AO22X1 U5106 ( .IN1(\read_value_mux[3][3] ), .IN2(n1643), .IN3(write_data[3]), .IN4(n3178), .Q(\words[3]/data_i[3] ) );
  AO22X1 U5107 ( .IN1(\read_value_mux[3][4] ), .IN2(n1643), .IN3(write_data[4]), .IN4(n3178), .Q(\words[3]/data_i[4] ) );
  AO22X1 U5108 ( .IN1(\read_value_mux[3][5] ), .IN2(n1643), .IN3(write_data[5]), .IN4(n3178), .Q(\words[3]/data_i[5] ) );
  AO22X1 U5109 ( .IN1(\read_value_mux[3][6] ), .IN2(n1643), .IN3(write_data[6]), .IN4(n3178), .Q(\words[3]/data_i[6] ) );
  AO22X1 U5110 ( .IN1(\read_value_mux[3][7] ), .IN2(n1643), .IN3(write_data[7]), .IN4(n3178), .Q(\words[3]/data_i[7] ) );
  AO22X1 U5111 ( .IN1(\read_value_mux[3][8] ), .IN2(n1643), .IN3(write_data[8]), .IN4(n3178), .Q(\words[3]/data_i[8] ) );
  AO22X1 U5112 ( .IN1(\read_value_mux[3][9] ), .IN2(n1643), .IN3(write_data[9]), .IN4(n3178), .Q(\words[3]/data_i[9] ) );
  AO21X1 U5113 ( .IN1(\words[3]/valid_o ), .IN2(n1743), .IN3(n3178), .Q(
        \words[3]/valid_i ) );
  AO22X1 U5114 ( .IN1(\read_value_mux[4][0] ), .IN2(n1634), .IN3(write_data[0]), .IN4(n3181), .Q(\words[4]/data_i[0] ) );
  AO22X1 U5115 ( .IN1(\read_value_mux[4][10] ), .IN2(n1634), .IN3(
        write_data[10]), .IN4(n3181), .Q(\words[4]/data_i[10] ) );
  AO22X1 U5116 ( .IN1(\read_value_mux[4][11] ), .IN2(n1634), .IN3(
        write_data[11]), .IN4(n3181), .Q(\words[4]/data_i[11] ) );
  AO22X1 U5117 ( .IN1(\read_value_mux[4][12] ), .IN2(n1634), .IN3(
        write_data[12]), .IN4(n3181), .Q(\words[4]/data_i[12] ) );
  AO22X1 U5118 ( .IN1(\read_value_mux[4][13] ), .IN2(n1634), .IN3(
        write_data[13]), .IN4(n3181), .Q(\words[4]/data_i[13] ) );
  AO22X1 U5119 ( .IN1(\read_value_mux[4][14] ), .IN2(n1634), .IN3(
        write_data[14]), .IN4(n3181), .Q(\words[4]/data_i[14] ) );
  AO22X1 U5120 ( .IN1(\read_value_mux[4][15] ), .IN2(n1634), .IN3(
        write_data[15]), .IN4(n3181), .Q(\words[4]/data_i[15] ) );
  AO22X1 U5121 ( .IN1(\read_value_mux[4][16] ), .IN2(n1634), .IN3(
        write_data[16]), .IN4(n3181), .Q(\words[4]/data_i[16] ) );
  AO22X1 U5122 ( .IN1(\read_value_mux[4][17] ), .IN2(n1634), .IN3(
        write_data[17]), .IN4(n3181), .Q(\words[4]/data_i[17] ) );
  AO22X1 U5123 ( .IN1(\read_value_mux[4][18] ), .IN2(n1634), .IN3(
        write_data[18]), .IN4(n3181), .Q(\words[4]/data_i[18] ) );
  AO22X1 U5124 ( .IN1(\read_value_mux[4][19] ), .IN2(n1634), .IN3(
        write_data[19]), .IN4(n3181), .Q(\words[4]/data_i[19] ) );
  AO22X1 U5125 ( .IN1(\read_value_mux[4][1] ), .IN2(n1634), .IN3(write_data[1]), .IN4(n3181), .Q(\words[4]/data_i[1] ) );
  AO22X1 U5126 ( .IN1(\read_value_mux[4][20] ), .IN2(n1634), .IN3(
        write_data[20]), .IN4(n3181), .Q(\words[4]/data_i[20] ) );
  AO22X1 U5127 ( .IN1(\read_value_mux[4][21] ), .IN2(n1634), .IN3(
        write_data[21]), .IN4(n3181), .Q(\words[4]/data_i[21] ) );
  AO22X1 U5128 ( .IN1(\read_value_mux[4][22] ), .IN2(n1634), .IN3(
        write_data[22]), .IN4(n3181), .Q(\words[4]/data_i[22] ) );
  AO22X1 U5129 ( .IN1(\read_value_mux[4][23] ), .IN2(n1634), .IN3(
        write_data[23]), .IN4(n3181), .Q(\words[4]/data_i[23] ) );
  AO22X1 U5130 ( .IN1(\read_value_mux[4][24] ), .IN2(n1634), .IN3(
        write_data[24]), .IN4(n3181), .Q(\words[4]/data_i[24] ) );
  AO22X1 U5131 ( .IN1(\read_value_mux[4][25] ), .IN2(n1634), .IN3(
        write_data[25]), .IN4(n3181), .Q(\words[4]/data_i[25] ) );
  AO22X1 U5132 ( .IN1(\read_value_mux[4][26] ), .IN2(n1634), .IN3(
        write_data[26]), .IN4(n3181), .Q(\words[4]/data_i[26] ) );
  AO22X1 U5133 ( .IN1(\read_value_mux[4][27] ), .IN2(n1634), .IN3(
        write_data[27]), .IN4(n3181), .Q(\words[4]/data_i[27] ) );
  AO22X1 U5134 ( .IN1(\read_value_mux[4][28] ), .IN2(n1634), .IN3(
        write_data[28]), .IN4(n3181), .Q(\words[4]/data_i[28] ) );
  AO22X1 U5135 ( .IN1(\read_value_mux[4][29] ), .IN2(n1634), .IN3(
        write_data[29]), .IN4(n3181), .Q(\words[4]/data_i[29] ) );
  AO22X1 U5136 ( .IN1(\read_value_mux[4][2] ), .IN2(n1634), .IN3(write_data[2]), .IN4(n3181), .Q(\words[4]/data_i[2] ) );
  AO22X1 U5137 ( .IN1(\read_value_mux[4][30] ), .IN2(n1634), .IN3(
        write_data[30]), .IN4(n3181), .Q(\words[4]/data_i[30] ) );
  AO22X1 U5138 ( .IN1(\read_value_mux[4][31] ), .IN2(n1634), .IN3(
        write_data[31]), .IN4(n3181), .Q(\words[4]/data_i[31] ) );
  AO22X1 U5139 ( .IN1(\read_value_mux[4][3] ), .IN2(n1634), .IN3(write_data[3]), .IN4(n3181), .Q(\words[4]/data_i[3] ) );
  AO22X1 U5140 ( .IN1(\read_value_mux[4][4] ), .IN2(n1634), .IN3(write_data[4]), .IN4(n3181), .Q(\words[4]/data_i[4] ) );
  AO22X1 U5141 ( .IN1(\read_value_mux[4][5] ), .IN2(n1634), .IN3(write_data[5]), .IN4(n3181), .Q(\words[4]/data_i[5] ) );
  AO22X1 U5142 ( .IN1(\read_value_mux[4][6] ), .IN2(n1634), .IN3(write_data[6]), .IN4(n3181), .Q(\words[4]/data_i[6] ) );
  AO22X1 U5143 ( .IN1(\read_value_mux[4][7] ), .IN2(n1634), .IN3(write_data[7]), .IN4(n3181), .Q(\words[4]/data_i[7] ) );
  AO22X1 U5144 ( .IN1(\read_value_mux[4][8] ), .IN2(n1634), .IN3(write_data[8]), .IN4(n3181), .Q(\words[4]/data_i[8] ) );
  AO22X1 U5145 ( .IN1(\read_value_mux[4][9] ), .IN2(n1634), .IN3(write_data[9]), .IN4(n3181), .Q(\words[4]/data_i[9] ) );
  AO21X1 U5146 ( .IN1(\words[4]/valid_o ), .IN2(n1743), .IN3(n3181), .Q(
        \words[4]/valid_i ) );
  AO22X1 U5147 ( .IN1(\read_value_mux[5][0] ), .IN2(n1616), .IN3(write_data[0]), .IN4(n3182), .Q(\words[5]/data_i[0] ) );
  AO22X1 U5148 ( .IN1(\read_value_mux[5][10] ), .IN2(n1616), .IN3(
        write_data[10]), .IN4(n3182), .Q(\words[5]/data_i[10] ) );
  AO22X1 U5149 ( .IN1(\read_value_mux[5][11] ), .IN2(n1616), .IN3(
        write_data[11]), .IN4(n3182), .Q(\words[5]/data_i[11] ) );
  AO22X1 U5150 ( .IN1(\read_value_mux[5][12] ), .IN2(n1616), .IN3(
        write_data[12]), .IN4(n3182), .Q(\words[5]/data_i[12] ) );
  AO22X1 U5151 ( .IN1(\read_value_mux[5][13] ), .IN2(n1616), .IN3(
        write_data[13]), .IN4(n3182), .Q(\words[5]/data_i[13] ) );
  AO22X1 U5152 ( .IN1(\read_value_mux[5][14] ), .IN2(n1616), .IN3(
        write_data[14]), .IN4(n3182), .Q(\words[5]/data_i[14] ) );
  AO22X1 U5153 ( .IN1(\read_value_mux[5][15] ), .IN2(n1616), .IN3(
        write_data[15]), .IN4(n3182), .Q(\words[5]/data_i[15] ) );
  AO22X1 U5154 ( .IN1(\read_value_mux[5][16] ), .IN2(n1616), .IN3(
        write_data[16]), .IN4(n3182), .Q(\words[5]/data_i[16] ) );
  AO22X1 U5155 ( .IN1(\read_value_mux[5][17] ), .IN2(n1616), .IN3(
        write_data[17]), .IN4(n3182), .Q(\words[5]/data_i[17] ) );
  AO22X1 U5156 ( .IN1(\read_value_mux[5][18] ), .IN2(n1616), .IN3(
        write_data[18]), .IN4(n3182), .Q(\words[5]/data_i[18] ) );
  AO22X1 U5157 ( .IN1(\read_value_mux[5][19] ), .IN2(n1616), .IN3(
        write_data[19]), .IN4(n3182), .Q(\words[5]/data_i[19] ) );
  AO22X1 U5158 ( .IN1(\read_value_mux[5][1] ), .IN2(n1616), .IN3(write_data[1]), .IN4(n3182), .Q(\words[5]/data_i[1] ) );
  AO22X1 U5159 ( .IN1(\read_value_mux[5][20] ), .IN2(n1616), .IN3(
        write_data[20]), .IN4(n3182), .Q(\words[5]/data_i[20] ) );
  AO22X1 U5160 ( .IN1(\read_value_mux[5][21] ), .IN2(n1616), .IN3(
        write_data[21]), .IN4(n3182), .Q(\words[5]/data_i[21] ) );
  AO22X1 U5161 ( .IN1(\read_value_mux[5][22] ), .IN2(n1616), .IN3(
        write_data[22]), .IN4(n3182), .Q(\words[5]/data_i[22] ) );
  AO22X1 U5162 ( .IN1(\read_value_mux[5][23] ), .IN2(n1616), .IN3(
        write_data[23]), .IN4(n3182), .Q(\words[5]/data_i[23] ) );
  AO22X1 U5163 ( .IN1(\read_value_mux[5][24] ), .IN2(n1616), .IN3(
        write_data[24]), .IN4(n3182), .Q(\words[5]/data_i[24] ) );
  AO22X1 U5164 ( .IN1(\read_value_mux[5][25] ), .IN2(n1616), .IN3(
        write_data[25]), .IN4(n3182), .Q(\words[5]/data_i[25] ) );
  AO22X1 U5165 ( .IN1(\read_value_mux[5][26] ), .IN2(n1616), .IN3(
        write_data[26]), .IN4(n3182), .Q(\words[5]/data_i[26] ) );
  AO22X1 U5166 ( .IN1(\read_value_mux[5][27] ), .IN2(n1616), .IN3(
        write_data[27]), .IN4(n3182), .Q(\words[5]/data_i[27] ) );
  AO22X1 U5167 ( .IN1(\read_value_mux[5][28] ), .IN2(n1616), .IN3(
        write_data[28]), .IN4(n3182), .Q(\words[5]/data_i[28] ) );
  AO22X1 U5168 ( .IN1(\read_value_mux[5][29] ), .IN2(n1616), .IN3(
        write_data[29]), .IN4(n3182), .Q(\words[5]/data_i[29] ) );
  AO22X1 U5169 ( .IN1(\read_value_mux[5][2] ), .IN2(n1616), .IN3(write_data[2]), .IN4(n3182), .Q(\words[5]/data_i[2] ) );
  AO22X1 U5170 ( .IN1(\read_value_mux[5][30] ), .IN2(n1616), .IN3(
        write_data[30]), .IN4(n3182), .Q(\words[5]/data_i[30] ) );
  AO22X1 U5171 ( .IN1(\read_value_mux[5][31] ), .IN2(n1616), .IN3(
        write_data[31]), .IN4(n3182), .Q(\words[5]/data_i[31] ) );
  AO22X1 U5172 ( .IN1(\read_value_mux[5][3] ), .IN2(n1616), .IN3(write_data[3]), .IN4(n3182), .Q(\words[5]/data_i[3] ) );
  AO22X1 U5173 ( .IN1(\read_value_mux[5][4] ), .IN2(n1616), .IN3(write_data[4]), .IN4(n3182), .Q(\words[5]/data_i[4] ) );
  AO22X1 U5174 ( .IN1(\read_value_mux[5][5] ), .IN2(n1616), .IN3(write_data[5]), .IN4(n3182), .Q(\words[5]/data_i[5] ) );
  AO22X1 U5175 ( .IN1(\read_value_mux[5][6] ), .IN2(n1616), .IN3(write_data[6]), .IN4(n3182), .Q(\words[5]/data_i[6] ) );
  AO22X1 U5176 ( .IN1(\read_value_mux[5][7] ), .IN2(n1616), .IN3(write_data[7]), .IN4(n3182), .Q(\words[5]/data_i[7] ) );
  AO22X1 U5177 ( .IN1(\read_value_mux[5][8] ), .IN2(n1616), .IN3(write_data[8]), .IN4(n3182), .Q(\words[5]/data_i[8] ) );
  AO22X1 U5178 ( .IN1(\read_value_mux[5][9] ), .IN2(n1616), .IN3(write_data[9]), .IN4(n3182), .Q(\words[5]/data_i[9] ) );
  AO21X1 U5179 ( .IN1(\words[5]/valid_o ), .IN2(n1743), .IN3(n3182), .Q(
        \words[5]/valid_i ) );
  AO22X1 U5180 ( .IN1(\read_value_mux[6][0] ), .IN2(n1644), .IN3(write_data[0]), .IN4(n3184), .Q(\words[6]/data_i[0] ) );
  AO22X1 U5181 ( .IN1(\read_value_mux[6][10] ), .IN2(n1644), .IN3(
        write_data[10]), .IN4(n3184), .Q(\words[6]/data_i[10] ) );
  AO22X1 U5182 ( .IN1(\read_value_mux[6][11] ), .IN2(n1644), .IN3(
        write_data[11]), .IN4(n3184), .Q(\words[6]/data_i[11] ) );
  AO22X1 U5183 ( .IN1(\read_value_mux[6][12] ), .IN2(n1644), .IN3(
        write_data[12]), .IN4(n3184), .Q(\words[6]/data_i[12] ) );
  AO22X1 U5184 ( .IN1(\read_value_mux[6][13] ), .IN2(n1644), .IN3(
        write_data[13]), .IN4(n3184), .Q(\words[6]/data_i[13] ) );
  AO22X1 U5185 ( .IN1(\read_value_mux[6][14] ), .IN2(n1644), .IN3(
        write_data[14]), .IN4(n3184), .Q(\words[6]/data_i[14] ) );
  AO22X1 U5186 ( .IN1(\read_value_mux[6][15] ), .IN2(n1644), .IN3(
        write_data[15]), .IN4(n3184), .Q(\words[6]/data_i[15] ) );
  AO22X1 U5187 ( .IN1(\read_value_mux[6][16] ), .IN2(n1644), .IN3(
        write_data[16]), .IN4(n3184), .Q(\words[6]/data_i[16] ) );
  AO22X1 U5188 ( .IN1(\read_value_mux[6][17] ), .IN2(n1644), .IN3(
        write_data[17]), .IN4(n3184), .Q(\words[6]/data_i[17] ) );
  AO22X1 U5189 ( .IN1(\read_value_mux[6][18] ), .IN2(n1644), .IN3(
        write_data[18]), .IN4(n3184), .Q(\words[6]/data_i[18] ) );
  AO22X1 U5190 ( .IN1(\read_value_mux[6][19] ), .IN2(n1644), .IN3(
        write_data[19]), .IN4(n3184), .Q(\words[6]/data_i[19] ) );
  AO22X1 U5191 ( .IN1(\read_value_mux[6][1] ), .IN2(n1644), .IN3(write_data[1]), .IN4(n3184), .Q(\words[6]/data_i[1] ) );
  AO22X1 U5192 ( .IN1(\read_value_mux[6][20] ), .IN2(n1644), .IN3(
        write_data[20]), .IN4(n3184), .Q(\words[6]/data_i[20] ) );
  AO22X1 U5193 ( .IN1(\read_value_mux[6][21] ), .IN2(n1644), .IN3(
        write_data[21]), .IN4(n3184), .Q(\words[6]/data_i[21] ) );
  AO22X1 U5194 ( .IN1(\read_value_mux[6][22] ), .IN2(n1644), .IN3(
        write_data[22]), .IN4(n3184), .Q(\words[6]/data_i[22] ) );
  AO22X1 U5195 ( .IN1(\read_value_mux[6][23] ), .IN2(n1644), .IN3(
        write_data[23]), .IN4(n3184), .Q(\words[6]/data_i[23] ) );
  AO22X1 U5196 ( .IN1(\read_value_mux[6][24] ), .IN2(n1644), .IN3(
        write_data[24]), .IN4(n3184), .Q(\words[6]/data_i[24] ) );
  AO22X1 U5197 ( .IN1(\read_value_mux[6][25] ), .IN2(n1644), .IN3(
        write_data[25]), .IN4(n3184), .Q(\words[6]/data_i[25] ) );
  AO22X1 U5198 ( .IN1(\read_value_mux[6][26] ), .IN2(n1644), .IN3(
        write_data[26]), .IN4(n3184), .Q(\words[6]/data_i[26] ) );
  AO22X1 U5199 ( .IN1(\read_value_mux[6][27] ), .IN2(n1644), .IN3(
        write_data[27]), .IN4(n3184), .Q(\words[6]/data_i[27] ) );
  AO22X1 U5200 ( .IN1(\read_value_mux[6][28] ), .IN2(n1644), .IN3(
        write_data[28]), .IN4(n3184), .Q(\words[6]/data_i[28] ) );
  AO22X1 U5201 ( .IN1(\read_value_mux[6][29] ), .IN2(n1644), .IN3(
        write_data[29]), .IN4(n3184), .Q(\words[6]/data_i[29] ) );
  AO22X1 U5202 ( .IN1(\read_value_mux[6][2] ), .IN2(n1644), .IN3(write_data[2]), .IN4(n3184), .Q(\words[6]/data_i[2] ) );
  AO22X1 U5203 ( .IN1(\read_value_mux[6][30] ), .IN2(n1644), .IN3(
        write_data[30]), .IN4(n3184), .Q(\words[6]/data_i[30] ) );
  AO22X1 U5204 ( .IN1(\read_value_mux[6][31] ), .IN2(n1644), .IN3(
        write_data[31]), .IN4(n3184), .Q(\words[6]/data_i[31] ) );
  AO22X1 U5205 ( .IN1(\read_value_mux[6][3] ), .IN2(n1644), .IN3(write_data[3]), .IN4(n3184), .Q(\words[6]/data_i[3] ) );
  AO22X1 U5206 ( .IN1(\read_value_mux[6][4] ), .IN2(n1644), .IN3(write_data[4]), .IN4(n3184), .Q(\words[6]/data_i[4] ) );
  AO22X1 U5207 ( .IN1(\read_value_mux[6][5] ), .IN2(n1644), .IN3(write_data[5]), .IN4(n3184), .Q(\words[6]/data_i[5] ) );
  AO22X1 U5208 ( .IN1(\read_value_mux[6][6] ), .IN2(n1644), .IN3(write_data[6]), .IN4(n3184), .Q(\words[6]/data_i[6] ) );
  AO22X1 U5209 ( .IN1(\read_value_mux[6][7] ), .IN2(n1644), .IN3(write_data[7]), .IN4(n3184), .Q(\words[6]/data_i[7] ) );
  AO22X1 U5210 ( .IN1(\read_value_mux[6][8] ), .IN2(n1644), .IN3(write_data[8]), .IN4(n3184), .Q(\words[6]/data_i[8] ) );
  AO22X1 U5211 ( .IN1(\read_value_mux[6][9] ), .IN2(n1644), .IN3(write_data[9]), .IN4(n3184), .Q(\words[6]/data_i[9] ) );
  AO21X1 U5212 ( .IN1(\words[6]/valid_o ), .IN2(n1743), .IN3(n3184), .Q(
        \words[6]/valid_i ) );
  AO22X1 U5213 ( .IN1(\read_value_mux[7][0] ), .IN2(n1645), .IN3(write_data[0]), .IN4(n3187), .Q(\words[7]/data_i[0] ) );
  AO22X1 U5214 ( .IN1(\read_value_mux[7][10] ), .IN2(n1645), .IN3(
        write_data[10]), .IN4(n3187), .Q(\words[7]/data_i[10] ) );
  AO22X1 U5215 ( .IN1(\read_value_mux[7][11] ), .IN2(n1645), .IN3(
        write_data[11]), .IN4(n3187), .Q(\words[7]/data_i[11] ) );
  AO22X1 U5216 ( .IN1(\read_value_mux[7][12] ), .IN2(n1645), .IN3(
        write_data[12]), .IN4(n3187), .Q(\words[7]/data_i[12] ) );
  AO22X1 U5217 ( .IN1(\read_value_mux[7][13] ), .IN2(n1645), .IN3(
        write_data[13]), .IN4(n3187), .Q(\words[7]/data_i[13] ) );
  AO22X1 U5218 ( .IN1(\read_value_mux[7][14] ), .IN2(n1645), .IN3(
        write_data[14]), .IN4(n3187), .Q(\words[7]/data_i[14] ) );
  AO22X1 U5219 ( .IN1(\read_value_mux[7][15] ), .IN2(n1645), .IN3(
        write_data[15]), .IN4(n3187), .Q(\words[7]/data_i[15] ) );
  AO22X1 U5220 ( .IN1(\read_value_mux[7][16] ), .IN2(n1645), .IN3(
        write_data[16]), .IN4(n3187), .Q(\words[7]/data_i[16] ) );
  AO22X1 U5221 ( .IN1(\read_value_mux[7][17] ), .IN2(n1645), .IN3(
        write_data[17]), .IN4(n3187), .Q(\words[7]/data_i[17] ) );
  AO22X1 U5222 ( .IN1(\read_value_mux[7][18] ), .IN2(n1645), .IN3(
        write_data[18]), .IN4(n3187), .Q(\words[7]/data_i[18] ) );
  AO22X1 U5223 ( .IN1(\read_value_mux[7][19] ), .IN2(n1645), .IN3(
        write_data[19]), .IN4(n3187), .Q(\words[7]/data_i[19] ) );
  AO22X1 U5224 ( .IN1(\read_value_mux[7][1] ), .IN2(n1645), .IN3(write_data[1]), .IN4(n3187), .Q(\words[7]/data_i[1] ) );
  AO22X1 U5225 ( .IN1(\read_value_mux[7][20] ), .IN2(n1645), .IN3(
        write_data[20]), .IN4(n3187), .Q(\words[7]/data_i[20] ) );
  AO22X1 U5226 ( .IN1(\read_value_mux[7][21] ), .IN2(n1645), .IN3(
        write_data[21]), .IN4(n3187), .Q(\words[7]/data_i[21] ) );
  AO22X1 U5227 ( .IN1(\read_value_mux[7][22] ), .IN2(n1645), .IN3(
        write_data[22]), .IN4(n3187), .Q(\words[7]/data_i[22] ) );
  AO22X1 U5228 ( .IN1(\read_value_mux[7][23] ), .IN2(n1645), .IN3(
        write_data[23]), .IN4(n3187), .Q(\words[7]/data_i[23] ) );
  AO22X1 U5229 ( .IN1(\read_value_mux[7][24] ), .IN2(n1645), .IN3(
        write_data[24]), .IN4(n3187), .Q(\words[7]/data_i[24] ) );
  AO22X1 U5230 ( .IN1(\read_value_mux[7][25] ), .IN2(n1645), .IN3(
        write_data[25]), .IN4(n3187), .Q(\words[7]/data_i[25] ) );
  AO22X1 U5231 ( .IN1(\read_value_mux[7][26] ), .IN2(n1645), .IN3(
        write_data[26]), .IN4(n3187), .Q(\words[7]/data_i[26] ) );
  AO22X1 U5232 ( .IN1(\read_value_mux[7][27] ), .IN2(n1645), .IN3(
        write_data[27]), .IN4(n3187), .Q(\words[7]/data_i[27] ) );
  AO22X1 U5233 ( .IN1(\read_value_mux[7][28] ), .IN2(n1645), .IN3(
        write_data[28]), .IN4(n3187), .Q(\words[7]/data_i[28] ) );
  AO22X1 U5234 ( .IN1(\read_value_mux[7][29] ), .IN2(n1645), .IN3(
        write_data[29]), .IN4(n3187), .Q(\words[7]/data_i[29] ) );
  AO22X1 U5235 ( .IN1(\read_value_mux[7][2] ), .IN2(n1645), .IN3(write_data[2]), .IN4(n3187), .Q(\words[7]/data_i[2] ) );
  AO22X1 U5236 ( .IN1(\read_value_mux[7][30] ), .IN2(n1645), .IN3(
        write_data[30]), .IN4(n3187), .Q(\words[7]/data_i[30] ) );
  AO22X1 U5237 ( .IN1(\read_value_mux[7][31] ), .IN2(n1645), .IN3(
        write_data[31]), .IN4(n3187), .Q(\words[7]/data_i[31] ) );
  AO22X1 U5238 ( .IN1(\read_value_mux[7][3] ), .IN2(n1645), .IN3(write_data[3]), .IN4(n3187), .Q(\words[7]/data_i[3] ) );
  AO22X1 U5239 ( .IN1(\read_value_mux[7][4] ), .IN2(n1645), .IN3(write_data[4]), .IN4(n3187), .Q(\words[7]/data_i[4] ) );
  AO22X1 U5240 ( .IN1(\read_value_mux[7][5] ), .IN2(n1645), .IN3(write_data[5]), .IN4(n3187), .Q(\words[7]/data_i[5] ) );
  AO22X1 U5241 ( .IN1(\read_value_mux[7][6] ), .IN2(n1645), .IN3(write_data[6]), .IN4(n3187), .Q(\words[7]/data_i[6] ) );
  AO22X1 U5242 ( .IN1(\read_value_mux[7][7] ), .IN2(n1645), .IN3(write_data[7]), .IN4(n3187), .Q(\words[7]/data_i[7] ) );
  AO22X1 U5243 ( .IN1(\read_value_mux[7][8] ), .IN2(n1645), .IN3(write_data[8]), .IN4(n3187), .Q(\words[7]/data_i[8] ) );
  AO22X1 U5244 ( .IN1(\read_value_mux[7][9] ), .IN2(n1645), .IN3(write_data[9]), .IN4(n3187), .Q(\words[7]/data_i[9] ) );
  AO21X1 U5245 ( .IN1(\words[7]/valid_o ), .IN2(n1743), .IN3(n3187), .Q(
        \words[7]/valid_i ) );
  AO22X1 U5246 ( .IN1(\read_value_mux[8][0] ), .IN2(n1635), .IN3(write_data[0]), .IN4(n3189), .Q(\words[8]/data_i[0] ) );
  AO22X1 U5247 ( .IN1(\read_value_mux[8][10] ), .IN2(n1635), .IN3(
        write_data[10]), .IN4(n3189), .Q(\words[8]/data_i[10] ) );
  AO22X1 U5248 ( .IN1(\read_value_mux[8][11] ), .IN2(n1635), .IN3(
        write_data[11]), .IN4(n3189), .Q(\words[8]/data_i[11] ) );
  AO22X1 U5249 ( .IN1(\read_value_mux[8][12] ), .IN2(n1635), .IN3(
        write_data[12]), .IN4(n3189), .Q(\words[8]/data_i[12] ) );
  AO22X1 U5250 ( .IN1(\read_value_mux[8][13] ), .IN2(n1635), .IN3(
        write_data[13]), .IN4(n3189), .Q(\words[8]/data_i[13] ) );
  AO22X1 U5251 ( .IN1(\read_value_mux[8][14] ), .IN2(n1635), .IN3(
        write_data[14]), .IN4(n3189), .Q(\words[8]/data_i[14] ) );
  AO22X1 U5252 ( .IN1(\read_value_mux[8][15] ), .IN2(n1635), .IN3(
        write_data[15]), .IN4(n3189), .Q(\words[8]/data_i[15] ) );
  AO22X1 U5253 ( .IN1(\read_value_mux[8][16] ), .IN2(n1635), .IN3(
        write_data[16]), .IN4(n3189), .Q(\words[8]/data_i[16] ) );
  AO22X1 U5254 ( .IN1(\read_value_mux[8][17] ), .IN2(n1635), .IN3(
        write_data[17]), .IN4(n3189), .Q(\words[8]/data_i[17] ) );
  AO22X1 U5255 ( .IN1(\read_value_mux[8][18] ), .IN2(n1635), .IN3(
        write_data[18]), .IN4(n3189), .Q(\words[8]/data_i[18] ) );
  AO22X1 U5256 ( .IN1(\read_value_mux[8][19] ), .IN2(n1635), .IN3(
        write_data[19]), .IN4(n3189), .Q(\words[8]/data_i[19] ) );
  AO22X1 U5257 ( .IN1(\read_value_mux[8][1] ), .IN2(n1635), .IN3(write_data[1]), .IN4(n3189), .Q(\words[8]/data_i[1] ) );
  AO22X1 U5258 ( .IN1(\read_value_mux[8][20] ), .IN2(n1635), .IN3(
        write_data[20]), .IN4(n3189), .Q(\words[8]/data_i[20] ) );
  AO22X1 U5259 ( .IN1(\read_value_mux[8][21] ), .IN2(n1635), .IN3(
        write_data[21]), .IN4(n3189), .Q(\words[8]/data_i[21] ) );
  AO22X1 U5260 ( .IN1(\read_value_mux[8][22] ), .IN2(n1635), .IN3(
        write_data[22]), .IN4(n3189), .Q(\words[8]/data_i[22] ) );
  AO22X1 U5261 ( .IN1(\read_value_mux[8][23] ), .IN2(n1635), .IN3(
        write_data[23]), .IN4(n3189), .Q(\words[8]/data_i[23] ) );
  AO22X1 U5262 ( .IN1(\read_value_mux[8][24] ), .IN2(n1635), .IN3(
        write_data[24]), .IN4(n3189), .Q(\words[8]/data_i[24] ) );
  AO22X1 U5263 ( .IN1(\read_value_mux[8][25] ), .IN2(n1635), .IN3(
        write_data[25]), .IN4(n3189), .Q(\words[8]/data_i[25] ) );
  AO22X1 U5264 ( .IN1(\read_value_mux[8][26] ), .IN2(n1635), .IN3(
        write_data[26]), .IN4(n3189), .Q(\words[8]/data_i[26] ) );
  AO22X1 U5265 ( .IN1(\read_value_mux[8][27] ), .IN2(n1635), .IN3(
        write_data[27]), .IN4(n3189), .Q(\words[8]/data_i[27] ) );
  AO22X1 U5266 ( .IN1(\read_value_mux[8][28] ), .IN2(n1635), .IN3(
        write_data[28]), .IN4(n3189), .Q(\words[8]/data_i[28] ) );
  AO22X1 U5267 ( .IN1(\read_value_mux[8][29] ), .IN2(n1635), .IN3(
        write_data[29]), .IN4(n3189), .Q(\words[8]/data_i[29] ) );
  AO22X1 U5268 ( .IN1(\read_value_mux[8][2] ), .IN2(n1635), .IN3(write_data[2]), .IN4(n3189), .Q(\words[8]/data_i[2] ) );
  AO22X1 U5269 ( .IN1(\read_value_mux[8][30] ), .IN2(n1635), .IN3(
        write_data[30]), .IN4(n3189), .Q(\words[8]/data_i[30] ) );
  AO22X1 U5270 ( .IN1(\read_value_mux[8][31] ), .IN2(n1635), .IN3(
        write_data[31]), .IN4(n3189), .Q(\words[8]/data_i[31] ) );
  AO22X1 U5271 ( .IN1(\read_value_mux[8][3] ), .IN2(n1635), .IN3(write_data[3]), .IN4(n3189), .Q(\words[8]/data_i[3] ) );
  AO22X1 U5272 ( .IN1(\read_value_mux[8][4] ), .IN2(n1635), .IN3(write_data[4]), .IN4(n3189), .Q(\words[8]/data_i[4] ) );
  AO22X1 U5273 ( .IN1(\read_value_mux[8][5] ), .IN2(n1635), .IN3(write_data[5]), .IN4(n3189), .Q(\words[8]/data_i[5] ) );
  AO22X1 U5274 ( .IN1(\read_value_mux[8][6] ), .IN2(n1635), .IN3(write_data[6]), .IN4(n3189), .Q(\words[8]/data_i[6] ) );
  AO22X1 U5275 ( .IN1(\read_value_mux[8][7] ), .IN2(n1635), .IN3(write_data[7]), .IN4(n3189), .Q(\words[8]/data_i[7] ) );
  AO22X1 U5276 ( .IN1(\read_value_mux[8][8] ), .IN2(n1635), .IN3(write_data[8]), .IN4(n3189), .Q(\words[8]/data_i[8] ) );
  AO22X1 U5277 ( .IN1(\read_value_mux[8][9] ), .IN2(n1635), .IN3(write_data[9]), .IN4(n3189), .Q(\words[8]/data_i[9] ) );
  AO21X1 U5278 ( .IN1(\words[8]/valid_o ), .IN2(n1743), .IN3(n3189), .Q(
        \words[8]/valid_i ) );
  AO22X1 U5279 ( .IN1(\read_value_mux[9][0] ), .IN2(n1636), .IN3(write_data[0]), .IN4(n3192), .Q(\words[9]/data_i[0] ) );
  AO22X1 U5280 ( .IN1(\read_value_mux[9][10] ), .IN2(n1636), .IN3(
        write_data[10]), .IN4(n3192), .Q(\words[9]/data_i[10] ) );
  AO22X1 U5281 ( .IN1(\read_value_mux[9][11] ), .IN2(n1636), .IN3(
        write_data[11]), .IN4(n3192), .Q(\words[9]/data_i[11] ) );
  AO22X1 U5282 ( .IN1(\read_value_mux[9][12] ), .IN2(n1636), .IN3(
        write_data[12]), .IN4(n3192), .Q(\words[9]/data_i[12] ) );
  AO22X1 U5283 ( .IN1(\read_value_mux[9][13] ), .IN2(n1636), .IN3(
        write_data[13]), .IN4(n3192), .Q(\words[9]/data_i[13] ) );
  AO22X1 U5284 ( .IN1(\read_value_mux[9][14] ), .IN2(n1636), .IN3(
        write_data[14]), .IN4(n3192), .Q(\words[9]/data_i[14] ) );
  AO22X1 U5285 ( .IN1(\read_value_mux[9][15] ), .IN2(n1636), .IN3(
        write_data[15]), .IN4(n3192), .Q(\words[9]/data_i[15] ) );
  AO22X1 U5286 ( .IN1(\read_value_mux[9][16] ), .IN2(n1636), .IN3(
        write_data[16]), .IN4(n3192), .Q(\words[9]/data_i[16] ) );
  AO22X1 U5287 ( .IN1(\read_value_mux[9][17] ), .IN2(n1636), .IN3(
        write_data[17]), .IN4(n3192), .Q(\words[9]/data_i[17] ) );
  AO22X1 U5288 ( .IN1(\read_value_mux[9][18] ), .IN2(n1636), .IN3(
        write_data[18]), .IN4(n3192), .Q(\words[9]/data_i[18] ) );
  AO22X1 U5289 ( .IN1(\read_value_mux[9][19] ), .IN2(n1636), .IN3(
        write_data[19]), .IN4(n3192), .Q(\words[9]/data_i[19] ) );
  AO22X1 U5290 ( .IN1(\read_value_mux[9][1] ), .IN2(n1636), .IN3(write_data[1]), .IN4(n3192), .Q(\words[9]/data_i[1] ) );
  AO22X1 U5291 ( .IN1(\read_value_mux[9][20] ), .IN2(n1636), .IN3(
        write_data[20]), .IN4(n3192), .Q(\words[9]/data_i[20] ) );
  AO22X1 U5292 ( .IN1(\read_value_mux[9][21] ), .IN2(n1636), .IN3(
        write_data[21]), .IN4(n3192), .Q(\words[9]/data_i[21] ) );
  AO22X1 U5293 ( .IN1(\read_value_mux[9][22] ), .IN2(n1636), .IN3(
        write_data[22]), .IN4(n3192), .Q(\words[9]/data_i[22] ) );
  AO22X1 U5294 ( .IN1(\read_value_mux[9][23] ), .IN2(n1636), .IN3(
        write_data[23]), .IN4(n3192), .Q(\words[9]/data_i[23] ) );
  AO22X1 U5295 ( .IN1(\read_value_mux[9][24] ), .IN2(n1636), .IN3(
        write_data[24]), .IN4(n3192), .Q(\words[9]/data_i[24] ) );
  AO22X1 U5296 ( .IN1(\read_value_mux[9][25] ), .IN2(n1636), .IN3(
        write_data[25]), .IN4(n3192), .Q(\words[9]/data_i[25] ) );
  AO22X1 U5297 ( .IN1(\read_value_mux[9][26] ), .IN2(n1636), .IN3(
        write_data[26]), .IN4(n3192), .Q(\words[9]/data_i[26] ) );
  AO22X1 U5298 ( .IN1(\read_value_mux[9][27] ), .IN2(n1636), .IN3(
        write_data[27]), .IN4(n3192), .Q(\words[9]/data_i[27] ) );
  AO22X1 U5299 ( .IN1(\read_value_mux[9][28] ), .IN2(n1636), .IN3(
        write_data[28]), .IN4(n3192), .Q(\words[9]/data_i[28] ) );
  AO22X1 U5300 ( .IN1(\read_value_mux[9][29] ), .IN2(n1636), .IN3(
        write_data[29]), .IN4(n3192), .Q(\words[9]/data_i[29] ) );
  AO22X1 U5301 ( .IN1(\read_value_mux[9][2] ), .IN2(n1636), .IN3(write_data[2]), .IN4(n3192), .Q(\words[9]/data_i[2] ) );
  AO22X1 U5302 ( .IN1(\read_value_mux[9][30] ), .IN2(n1636), .IN3(
        write_data[30]), .IN4(n3192), .Q(\words[9]/data_i[30] ) );
  AO22X1 U5303 ( .IN1(\read_value_mux[9][31] ), .IN2(n1636), .IN3(
        write_data[31]), .IN4(n3192), .Q(\words[9]/data_i[31] ) );
  AO22X1 U5304 ( .IN1(\read_value_mux[9][3] ), .IN2(n1636), .IN3(write_data[3]), .IN4(n3192), .Q(\words[9]/data_i[3] ) );
  AO22X1 U5305 ( .IN1(\read_value_mux[9][4] ), .IN2(n1636), .IN3(write_data[4]), .IN4(n3192), .Q(\words[9]/data_i[4] ) );
  AO22X1 U5306 ( .IN1(\read_value_mux[9][5] ), .IN2(n1636), .IN3(write_data[5]), .IN4(n3192), .Q(\words[9]/data_i[5] ) );
  AO22X1 U5307 ( .IN1(\read_value_mux[9][6] ), .IN2(n1636), .IN3(write_data[6]), .IN4(n3192), .Q(\words[9]/data_i[6] ) );
  AO22X1 U5308 ( .IN1(\read_value_mux[9][7] ), .IN2(n1636), .IN3(write_data[7]), .IN4(n3192), .Q(\words[9]/data_i[7] ) );
  AO22X1 U5309 ( .IN1(\read_value_mux[9][8] ), .IN2(n1636), .IN3(write_data[8]), .IN4(n3192), .Q(\words[9]/data_i[8] ) );
  AO22X1 U5310 ( .IN1(\read_value_mux[9][9] ), .IN2(n1636), .IN3(write_data[9]), .IN4(n3192), .Q(\words[9]/data_i[9] ) );
  AO21X1 U5311 ( .IN1(\words[9]/valid_o ), .IN2(n1743), .IN3(n3192), .Q(
        \words[9]/valid_i ) );
endmodule

