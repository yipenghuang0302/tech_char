
module cam_word_0 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  OAI22D0 U3 ( .A1(n46), .A2(search_data[19]), .B1(n47), .B2(search_data[22]), 
        .ZN(n1) );
  AOI221D0 U4 ( .A1(n46), .A2(search_data[19]), .B1(search_data[22]), .B2(n47), 
        .C(n1), .ZN(n2) );
  CKND0 U5 ( .I(read_value[21]), .ZN(n3) );
  CKND0 U6 ( .I(read_value[8]), .ZN(n4) );
  OAI22D0 U7 ( .A1(search_data[21]), .A2(n3), .B1(search_data[8]), .B2(n4), 
        .ZN(n5) );
  AOI221D0 U8 ( .A1(n4), .A2(search_data[8]), .B1(n3), .B2(search_data[21]), 
        .C(n5), .ZN(n6) );
  OAI22D0 U9 ( .A1(n50), .A2(search_data[15]), .B1(n51), .B2(search_data[18]), 
        .ZN(n7) );
  AOI221D0 U10 ( .A1(n50), .A2(search_data[15]), .B1(search_data[18]), .B2(n51), .C(n7), .ZN(n8) );
  OAI22D0 U11 ( .A1(n48), .A2(search_data[17]), .B1(n49), .B2(search_data[20]), 
        .ZN(n9) );
  AOI221D0 U12 ( .A1(n48), .A2(search_data[17]), .B1(search_data[20]), .B2(n49), .C(n9), .ZN(n10) );
  ND4D0 U13 ( .A1(n2), .A2(n6), .A3(n8), .A4(n10), .ZN(n11) );
  CKND0 U14 ( .I(read_value[27]), .ZN(n12) );
  CKND0 U15 ( .I(read_value[30]), .ZN(n13) );
  OAI22D0 U16 ( .A1(search_data[27]), .A2(n12), .B1(search_data[30]), .B2(n13), 
        .ZN(n14) );
  AOI221D0 U17 ( .A1(n13), .A2(search_data[30]), .B1(n12), .B2(search_data[27]), .C(n14), .ZN(n15) );
  CKND0 U18 ( .I(read_value[29]), .ZN(n16) );
  CKND0 U19 ( .I(read_value[31]), .ZN(n17) );
  OAI22D0 U20 ( .A1(search_data[29]), .A2(n16), .B1(search_data[31]), .B2(n17), 
        .ZN(n18) );
  AOI221D0 U21 ( .A1(n17), .A2(search_data[31]), .B1(n16), .B2(search_data[29]), .C(n18), .ZN(n19) );
  CKND0 U22 ( .I(read_value[23]), .ZN(n20) );
  CKND0 U23 ( .I(read_value[26]), .ZN(n21) );
  OAI22D0 U24 ( .A1(search_data[23]), .A2(n20), .B1(search_data[26]), .B2(n21), 
        .ZN(n22) );
  AOI221D0 U25 ( .A1(n21), .A2(search_data[26]), .B1(n20), .B2(search_data[23]), .C(n22), .ZN(n23) );
  CKND0 U26 ( .I(read_value[24]), .ZN(n24) );
  CKND0 U27 ( .I(read_value[28]), .ZN(n25) );
  OAI22D0 U28 ( .A1(search_data[24]), .A2(n24), .B1(search_data[28]), .B2(n25), 
        .ZN(n26) );
  AOI221D0 U29 ( .A1(n25), .A2(search_data[28]), .B1(n24), .B2(search_data[24]), .C(n26), .ZN(n27) );
  ND4D0 U30 ( .A1(n15), .A2(n19), .A3(n23), .A4(n27), .ZN(n28) );
  OAI22D0 U31 ( .A1(n60), .A2(search_data[5]), .B1(n61), .B2(search_data[7]), 
        .ZN(n29) );
  AOI221D0 U32 ( .A1(n60), .A2(search_data[5]), .B1(search_data[7]), .B2(n61), 
        .C(n29), .ZN(n30) );
  OAI22D0 U33 ( .A1(n62), .A2(search_data[2]), .B1(n63), .B2(search_data[16]), 
        .ZN(n31) );
  AOI221D0 U34 ( .A1(n62), .A2(search_data[2]), .B1(search_data[16]), .B2(n63), 
        .C(n31), .ZN(n32) );
  OA22D0 U35 ( .A1(search_data[3]), .A2(n66), .B1(search_data[6]), .B2(n65), 
        .Z(n33) );
  OA22D0 U36 ( .A1(search_data[1]), .A2(n69), .B1(search_data[4]), .B2(n68), 
        .Z(n34) );
  AN4D0 U37 ( .A1(n64), .A2(n33), .A3(n67), .A4(n34), .Z(n35) );
  ND4D0 U38 ( .A1(n30), .A2(search), .A3(n32), .A4(n35), .ZN(n36) );
  OAI22D0 U39 ( .A1(n54), .A2(search_data[11]), .B1(n55), .B2(search_data[14]), 
        .ZN(n37) );
  AOI221D0 U40 ( .A1(n54), .A2(search_data[11]), .B1(search_data[14]), .B2(n55), .C(n37), .ZN(n38) );
  OAI22D0 U41 ( .A1(n52), .A2(search_data[13]), .B1(n53), .B2(search_data[0]), 
        .ZN(n39) );
  AOI221D0 U42 ( .A1(n52), .A2(search_data[13]), .B1(search_data[0]), .B2(n53), 
        .C(n39), .ZN(n40) );
  OAI22D0 U43 ( .A1(n58), .A2(search_data[25]), .B1(n59), .B2(search_data[10]), 
        .ZN(n41) );
  AOI221D0 U44 ( .A1(n58), .A2(search_data[25]), .B1(search_data[10]), .B2(n59), .C(n41), .ZN(n42) );
  OAI22D0 U45 ( .A1(n56), .A2(search_data[9]), .B1(n57), .B2(search_data[12]), 
        .ZN(n43) );
  AOI221D0 U46 ( .A1(n56), .A2(search_data[9]), .B1(search_data[12]), .B2(n57), 
        .C(n43), .ZN(n44) );
  ND4D0 U47 ( .A1(n38), .A2(n40), .A3(n42), .A4(n44), .ZN(n45) );
  NR4D0 U48 ( .A1(n11), .A2(n28), .A3(n36), .A4(n45), .ZN(search_results) );
  AN3D0 U49 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results)
         );
  AO21D0 U50 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U51 ( .A1(reset), .A2(n70), .ZN(n71) );
  AOI21D2 U52 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  CKND2D1 U53 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  CKND0 U54 ( .I(read_value[3]), .ZN(n66) );
  CKND1 U55 ( .I(read_value[22]), .ZN(n47) );
  CKND1 U56 ( .I(read_value[25]), .ZN(n58) );
  CKND1 U57 ( .I(read_value[19]), .ZN(n46) );
  CKND0 U58 ( .I(read_value[6]), .ZN(n65) );
  CKND1 U59 ( .I(read_value[16]), .ZN(n63) );
  CKND1 U60 ( .I(read_value[5]), .ZN(n60) );
  CKND1 U61 ( .I(read_value[7]), .ZN(n61) );
  CKND1 U62 ( .I(read_value[2]), .ZN(n62) );
  CKND1 U63 ( .I(read_value[12]), .ZN(n57) );
  CKND1 U64 ( .I(read_value[0]), .ZN(n53) );
  CKND1 U65 ( .I(read_value[13]), .ZN(n52) );
  CKND1 U66 ( .I(read_value[15]), .ZN(n50) );
  CKND1 U67 ( .I(read_value[14]), .ZN(n55) );
  CKND1 U68 ( .I(read_value[11]), .ZN(n54) );
  CKND1 U69 ( .I(read_value[10]), .ZN(n59) );
  CKND0 U70 ( .I(read_value[1]), .ZN(n69) );
  CKND1 U71 ( .I(read_value[20]), .ZN(n49) );
  CKND1 U72 ( .I(read_value[17]), .ZN(n48) );
  CKND0 U73 ( .I(read_value[4]), .ZN(n68) );
  CKND1 U74 ( .I(read_value[18]), .ZN(n51) );
  CKND1 U75 ( .I(read_value[9]), .ZN(n56) );
  AO22D0 U76 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U77 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U78 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U79 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U80 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U81 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U82 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U83 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U84 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U85 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U86 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U87 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U88 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U89 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U90 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U91 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U92 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U93 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U94 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U95 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AOI22D1 U96 ( .A1(search_data[1]), .A2(n69), .B1(search_data[4]), .B2(n68), 
        .ZN(n67) );
  AOI22D1 U97 ( .A1(search_data[3]), .A2(n66), .B1(search_data[6]), .B2(n65), 
        .ZN(n64) );
  AO22D0 U98 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U99 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U100 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), 
        .Z(data_i[2]) );
  AO22D0 U101 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), 
        .Z(data_i[3]) );
  AO22D0 U102 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), 
        .Z(data_i[4]) );
  AO22D0 U103 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), 
        .Z(data_i[5]) );
  AO22D0 U104 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), 
        .Z(data_i[6]) );
  AO22D0 U105 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U106 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U107 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U108 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_1 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AOI221D0 U4 ( .A1(n9), .A2(search_data[31]), .B1(search_data[29]), .B2(n8), 
        .C(n7), .ZN(n22) );
  AOI221D0 U5 ( .A1(n12), .A2(search_data[30]), .B1(search_data[27]), .B2(n11), 
        .C(n10), .ZN(n21) );
  AOI221D0 U6 ( .A1(n15), .A2(search_data[28]), .B1(search_data[24]), .B2(n14), 
        .C(n13), .ZN(n20) );
  AOI221D0 U7 ( .A1(n18), .A2(search_data[26]), .B1(search_data[23]), .B2(n17), 
        .C(n16), .ZN(n19) );
  AOI221D0 U8 ( .A1(n25), .A2(search_data[8]), .B1(search_data[21]), .B2(n24), 
        .C(n23), .ZN(n38) );
  AOI221D0 U9 ( .A1(n28), .A2(search_data[22]), .B1(search_data[19]), .B2(n27), 
        .C(n26), .ZN(n37) );
  AOI221D0 U10 ( .A1(n31), .A2(search_data[20]), .B1(search_data[17]), .B2(n30), .C(n29), .ZN(n36) );
  AOI221D0 U11 ( .A1(n34), .A2(search_data[18]), .B1(search_data[15]), .B2(n33), .C(n32), .ZN(n35) );
  AOI221D0 U12 ( .A1(n41), .A2(search_data[0]), .B1(search_data[13]), .B2(n40), 
        .C(n39), .ZN(n54) );
  AOI221D0 U13 ( .A1(n44), .A2(search_data[14]), .B1(search_data[11]), .B2(n43), .C(n42), .ZN(n53) );
  AOI221D0 U14 ( .A1(n47), .A2(search_data[12]), .B1(search_data[9]), .B2(n46), 
        .C(n45), .ZN(n52) );
  AOI221D0 U15 ( .A1(n50), .A2(search_data[10]), .B1(search_data[25]), .B2(n49), .C(n48), .ZN(n51) );
  AOI221D0 U16 ( .A1(n57), .A2(search_data[7]), .B1(search_data[5]), .B2(n56), 
        .C(n55), .ZN(n65) );
  AOI221D0 U17 ( .A1(n60), .A2(search_data[16]), .B1(search_data[2]), .B2(n59), 
        .C(n58), .ZN(n64) );
  CKND0 U18 ( .I(read_value[4]), .ZN(n1) );
  CKND0 U19 ( .I(read_value[1]), .ZN(n2) );
  AOI22D0 U20 ( .A1(search_data[4]), .A2(n1), .B1(search_data[1]), .B2(n2), 
        .ZN(n3) );
  OAI221D0 U21 ( .A1(n1), .A2(search_data[4]), .B1(n2), .B2(search_data[1]), 
        .C(n3), .ZN(n61) );
  CKND0 U22 ( .I(read_value[6]), .ZN(n4) );
  CKND0 U23 ( .I(read_value[3]), .ZN(n5) );
  AOI22D0 U24 ( .A1(search_data[6]), .A2(n4), .B1(search_data[3]), .B2(n5), 
        .ZN(n6) );
  OAI221D0 U25 ( .A1(n4), .A2(search_data[6]), .B1(n5), .B2(search_data[3]), 
        .C(n6), .ZN(n62) );
  AN3D0 U26 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results)
         );
  AO21D0 U27 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U28 ( .A1(reset), .A2(n70), .ZN(n71) );
  CKND2D1 U29 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  AOI21D2 U30 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  CKND0 U31 ( .I(read_value[27]), .ZN(n11) );
  CKND0 U32 ( .I(read_value[30]), .ZN(n12) );
  CKND0 U33 ( .I(read_value[29]), .ZN(n8) );
  CKND0 U34 ( .I(read_value[31]), .ZN(n9) );
  CKND0 U35 ( .I(read_value[15]), .ZN(n33) );
  CKND0 U36 ( .I(read_value[18]), .ZN(n34) );
  CKND0 U37 ( .I(read_value[17]), .ZN(n30) );
  CKND0 U38 ( .I(read_value[20]), .ZN(n31) );
  CKND0 U39 ( .I(read_value[19]), .ZN(n27) );
  CKND0 U40 ( .I(read_value[22]), .ZN(n28) );
  CKND0 U41 ( .I(read_value[21]), .ZN(n24) );
  CKND0 U42 ( .I(read_value[8]), .ZN(n25) );
  CKND0 U43 ( .I(read_value[23]), .ZN(n17) );
  CKND0 U44 ( .I(read_value[26]), .ZN(n18) );
  CKND0 U45 ( .I(read_value[24]), .ZN(n14) );
  CKND0 U46 ( .I(read_value[28]), .ZN(n15) );
  CKND0 U47 ( .I(read_value[10]), .ZN(n50) );
  CKND0 U48 ( .I(read_value[25]), .ZN(n49) );
  CKND0 U49 ( .I(read_value[7]), .ZN(n57) );
  CKND0 U50 ( .I(read_value[5]), .ZN(n56) );
  CKND0 U51 ( .I(read_value[16]), .ZN(n60) );
  CKND0 U52 ( .I(read_value[2]), .ZN(n59) );
  CKND0 U53 ( .I(read_value[14]), .ZN(n44) );
  CKND0 U54 ( .I(read_value[11]), .ZN(n43) );
  CKND0 U55 ( .I(read_value[13]), .ZN(n40) );
  CKND0 U56 ( .I(read_value[12]), .ZN(n47) );
  CKND0 U57 ( .I(read_value[0]), .ZN(n41) );
  CKND0 U58 ( .I(read_value[9]), .ZN(n46) );
  AO22D0 U59 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U60 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U61 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U62 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U63 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U64 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U65 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U66 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U67 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U68 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U69 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U70 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U71 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U72 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U73 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U74 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U75 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U76 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U77 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U78 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  ND4D1 U79 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  NR2D1 U80 ( .A1(n62), .A2(n61), .ZN(n63) );
  OAI22D1 U81 ( .A1(n60), .A2(search_data[16]), .B1(n59), .B2(search_data[2]), 
        .ZN(n58) );
  OAI22D1 U82 ( .A1(n57), .A2(search_data[7]), .B1(n56), .B2(search_data[5]), 
        .ZN(n55) );
  ND4D1 U83 ( .A1(n54), .A2(n53), .A3(n52), .A4(n51), .ZN(n67) );
  OAI22D1 U84 ( .A1(n50), .A2(search_data[10]), .B1(n49), .B2(search_data[25]), 
        .ZN(n48) );
  OAI22D1 U85 ( .A1(n47), .A2(search_data[12]), .B1(n46), .B2(search_data[9]), 
        .ZN(n45) );
  OAI22D1 U86 ( .A1(n44), .A2(search_data[14]), .B1(n43), .B2(search_data[11]), 
        .ZN(n42) );
  OAI22D1 U87 ( .A1(n41), .A2(search_data[0]), .B1(n40), .B2(search_data[13]), 
        .ZN(n39) );
  ND4D1 U88 ( .A1(n38), .A2(n37), .A3(n36), .A4(n35), .ZN(n68) );
  OAI22D1 U89 ( .A1(n34), .A2(search_data[18]), .B1(n33), .B2(search_data[15]), 
        .ZN(n32) );
  OAI22D1 U90 ( .A1(n31), .A2(search_data[20]), .B1(n30), .B2(search_data[17]), 
        .ZN(n29) );
  OAI22D1 U91 ( .A1(n28), .A2(search_data[22]), .B1(n27), .B2(search_data[19]), 
        .ZN(n26) );
  OAI22D1 U92 ( .A1(n25), .A2(search_data[8]), .B1(n24), .B2(search_data[21]), 
        .ZN(n23) );
  ND4D1 U93 ( .A1(n22), .A2(n21), .A3(n20), .A4(n19), .ZN(n69) );
  OAI22D1 U94 ( .A1(n18), .A2(search_data[26]), .B1(n17), .B2(search_data[23]), 
        .ZN(n16) );
  OAI22D1 U95 ( .A1(n15), .A2(search_data[28]), .B1(n14), .B2(search_data[24]), 
        .ZN(n13) );
  OAI22D1 U96 ( .A1(n12), .A2(search_data[30]), .B1(n11), .B2(search_data[27]), 
        .ZN(n10) );
  OAI22D1 U97 ( .A1(n9), .A2(search_data[31]), .B1(n8), .B2(search_data[29]), 
        .ZN(n7) );
  AO22D0 U98 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U99 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U100 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), 
        .Z(data_i[2]) );
  AO22D0 U101 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), 
        .Z(data_i[3]) );
  AO22D0 U102 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), 
        .Z(data_i[4]) );
  AO22D0 U103 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), 
        .Z(data_i[5]) );
  AO22D0 U104 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), 
        .Z(data_i[6]) );
  AO22D0 U105 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U106 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U107 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U108 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_2 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AOI221D0 U4 ( .A1(n3), .A2(search_data[31]), .B1(search_data[29]), .B2(n2), 
        .C(n1), .ZN(n16) );
  AOI221D0 U5 ( .A1(n6), .A2(search_data[30]), .B1(search_data[27]), .B2(n5), 
        .C(n4), .ZN(n15) );
  AOI221D0 U6 ( .A1(n9), .A2(search_data[28]), .B1(search_data[24]), .B2(n8), 
        .C(n7), .ZN(n14) );
  AOI221D0 U7 ( .A1(n12), .A2(search_data[26]), .B1(search_data[23]), .B2(n11), 
        .C(n10), .ZN(n13) );
  AOI221D0 U8 ( .A1(n19), .A2(search_data[8]), .B1(search_data[21]), .B2(n18), 
        .C(n17), .ZN(n32) );
  AOI221D0 U9 ( .A1(n22), .A2(search_data[22]), .B1(search_data[19]), .B2(n21), 
        .C(n20), .ZN(n31) );
  AOI221D0 U10 ( .A1(n25), .A2(search_data[20]), .B1(search_data[17]), .B2(n24), .C(n23), .ZN(n30) );
  AOI221D0 U11 ( .A1(n28), .A2(search_data[18]), .B1(search_data[15]), .B2(n27), .C(n26), .ZN(n29) );
  AOI221D0 U12 ( .A1(n35), .A2(search_data[0]), .B1(search_data[13]), .B2(n34), 
        .C(n33), .ZN(n48) );
  AOI221D0 U13 ( .A1(n38), .A2(search_data[14]), .B1(search_data[11]), .B2(n37), .C(n36), .ZN(n47) );
  AOI221D0 U14 ( .A1(n41), .A2(search_data[12]), .B1(search_data[9]), .B2(n40), 
        .C(n39), .ZN(n46) );
  AOI221D0 U15 ( .A1(n44), .A2(search_data[10]), .B1(search_data[25]), .B2(n43), .C(n42), .ZN(n45) );
  AOI221D0 U16 ( .A1(n51), .A2(search_data[7]), .B1(search_data[5]), .B2(n50), 
        .C(n49), .ZN(n65) );
  AOI221D0 U17 ( .A1(n54), .A2(search_data[16]), .B1(search_data[2]), .B2(n53), 
        .C(n52), .ZN(n64) );
  OAI221D0 U18 ( .A1(n57), .A2(search_data[3]), .B1(n56), .B2(search_data[6]), 
        .C(n55), .ZN(n62) );
  OAI221D0 U19 ( .A1(n60), .A2(search_data[1]), .B1(n59), .B2(search_data[4]), 
        .C(n58), .ZN(n61) );
  AN3D0 U20 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results)
         );
  AO21D0 U21 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U22 ( .A1(reset), .A2(n70), .ZN(n71) );
  CKND2D1 U23 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  AOI21D2 U24 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  CKND0 U25 ( .I(read_value[8]), .ZN(n19) );
  CKND0 U26 ( .I(read_value[21]), .ZN(n18) );
  CKND0 U27 ( .I(read_value[30]), .ZN(n6) );
  CKND0 U28 ( .I(read_value[22]), .ZN(n22) );
  CKND0 U29 ( .I(read_value[12]), .ZN(n41) );
  CKND0 U30 ( .I(read_value[24]), .ZN(n8) );
  CKND0 U31 ( .I(read_value[31]), .ZN(n3) );
  CKND0 U32 ( .I(read_value[26]), .ZN(n12) );
  CKND0 U33 ( .I(read_value[23]), .ZN(n11) );
  CKND0 U34 ( .I(read_value[29]), .ZN(n2) );
  CKND0 U35 ( .I(read_value[28]), .ZN(n9) );
  CKND0 U36 ( .I(read_value[19]), .ZN(n21) );
  CKND0 U37 ( .I(read_value[1]), .ZN(n60) );
  CKND0 U38 ( .I(read_value[6]), .ZN(n56) );
  CKND0 U39 ( .I(read_value[0]), .ZN(n35) );
  CKND0 U40 ( .I(read_value[3]), .ZN(n57) );
  CKND0 U41 ( .I(read_value[13]), .ZN(n34) );
  CKND0 U42 ( .I(read_value[2]), .ZN(n53) );
  CKND0 U43 ( .I(read_value[16]), .ZN(n54) );
  CKND0 U44 ( .I(read_value[5]), .ZN(n50) );
  CKND0 U45 ( .I(read_value[14]), .ZN(n38) );
  CKND0 U46 ( .I(read_value[7]), .ZN(n51) );
  CKND0 U47 ( .I(read_value[11]), .ZN(n37) );
  CKND0 U48 ( .I(read_value[25]), .ZN(n43) );
  CKND0 U49 ( .I(read_value[10]), .ZN(n44) );
  CKND0 U50 ( .I(read_value[9]), .ZN(n40) );
  CKND0 U51 ( .I(read_value[20]), .ZN(n25) );
  CKND0 U52 ( .I(read_value[17]), .ZN(n24) );
  CKND0 U53 ( .I(read_value[27]), .ZN(n5) );
  CKND0 U54 ( .I(read_value[18]), .ZN(n28) );
  CKND0 U55 ( .I(read_value[15]), .ZN(n27) );
  CKND0 U56 ( .I(read_value[4]), .ZN(n59) );
  AO22D0 U57 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U58 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U59 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U60 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U61 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U62 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U63 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U64 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U65 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U66 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U67 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U68 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U69 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U70 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U71 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U72 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U73 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U74 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U75 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U76 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  ND4D1 U77 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  NR2D1 U78 ( .A1(n62), .A2(n61), .ZN(n63) );
  AOI22D1 U79 ( .A1(search_data[1]), .A2(n60), .B1(search_data[4]), .B2(n59), 
        .ZN(n58) );
  AOI22D1 U80 ( .A1(search_data[3]), .A2(n57), .B1(search_data[6]), .B2(n56), 
        .ZN(n55) );
  OAI22D1 U81 ( .A1(n54), .A2(search_data[16]), .B1(n53), .B2(search_data[2]), 
        .ZN(n52) );
  OAI22D1 U82 ( .A1(n51), .A2(search_data[7]), .B1(n50), .B2(search_data[5]), 
        .ZN(n49) );
  ND4D1 U83 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .ZN(n67) );
  OAI22D1 U84 ( .A1(n44), .A2(search_data[10]), .B1(n43), .B2(search_data[25]), 
        .ZN(n42) );
  OAI22D1 U85 ( .A1(n41), .A2(search_data[12]), .B1(n40), .B2(search_data[9]), 
        .ZN(n39) );
  OAI22D1 U86 ( .A1(n38), .A2(search_data[14]), .B1(n37), .B2(search_data[11]), 
        .ZN(n36) );
  OAI22D1 U87 ( .A1(n35), .A2(search_data[0]), .B1(n34), .B2(search_data[13]), 
        .ZN(n33) );
  ND4D1 U88 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .ZN(n68) );
  OAI22D1 U89 ( .A1(n28), .A2(search_data[18]), .B1(n27), .B2(search_data[15]), 
        .ZN(n26) );
  OAI22D1 U90 ( .A1(n25), .A2(search_data[20]), .B1(n24), .B2(search_data[17]), 
        .ZN(n23) );
  OAI22D1 U91 ( .A1(n22), .A2(search_data[22]), .B1(n21), .B2(search_data[19]), 
        .ZN(n20) );
  OAI22D1 U92 ( .A1(n19), .A2(search_data[8]), .B1(n18), .B2(search_data[21]), 
        .ZN(n17) );
  ND4D1 U93 ( .A1(n16), .A2(n15), .A3(n14), .A4(n13), .ZN(n69) );
  OAI22D1 U94 ( .A1(n12), .A2(search_data[26]), .B1(n11), .B2(search_data[23]), 
        .ZN(n10) );
  OAI22D1 U95 ( .A1(n9), .A2(search_data[28]), .B1(n8), .B2(search_data[24]), 
        .ZN(n7) );
  OAI22D1 U96 ( .A1(n6), .A2(search_data[30]), .B1(n5), .B2(search_data[27]), 
        .ZN(n4) );
  OAI22D1 U97 ( .A1(n3), .A2(search_data[31]), .B1(n2), .B2(search_data[29]), 
        .ZN(n1) );
  AO22D0 U98 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U99 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U100 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), 
        .Z(data_i[2]) );
  AO22D0 U101 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), 
        .Z(data_i[3]) );
  AO22D0 U102 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), 
        .Z(data_i[4]) );
  AO22D0 U103 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), 
        .Z(data_i[5]) );
  AO22D0 U104 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), 
        .Z(data_i[6]) );
  AO22D0 U105 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U106 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U107 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U108 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_3 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AOI221D0 U4 ( .A1(n3), .A2(search_data[31]), .B1(search_data[29]), .B2(n2), 
        .C(n1), .ZN(n16) );
  AOI221D0 U5 ( .A1(n6), .A2(search_data[30]), .B1(search_data[27]), .B2(n5), 
        .C(n4), .ZN(n15) );
  AOI221D0 U6 ( .A1(n9), .A2(search_data[28]), .B1(search_data[24]), .B2(n8), 
        .C(n7), .ZN(n14) );
  AOI221D0 U7 ( .A1(n12), .A2(search_data[26]), .B1(search_data[23]), .B2(n11), 
        .C(n10), .ZN(n13) );
  AOI221D0 U8 ( .A1(n19), .A2(search_data[8]), .B1(search_data[21]), .B2(n18), 
        .C(n17), .ZN(n32) );
  AOI221D0 U9 ( .A1(n22), .A2(search_data[22]), .B1(search_data[19]), .B2(n21), 
        .C(n20), .ZN(n31) );
  AOI221D0 U10 ( .A1(n25), .A2(search_data[20]), .B1(search_data[17]), .B2(n24), .C(n23), .ZN(n30) );
  AOI221D0 U11 ( .A1(n28), .A2(search_data[18]), .B1(search_data[15]), .B2(n27), .C(n26), .ZN(n29) );
  AOI221D0 U12 ( .A1(n35), .A2(search_data[0]), .B1(search_data[13]), .B2(n34), 
        .C(n33), .ZN(n48) );
  AOI221D0 U13 ( .A1(n38), .A2(search_data[14]), .B1(search_data[11]), .B2(n37), .C(n36), .ZN(n47) );
  AOI221D0 U14 ( .A1(n41), .A2(search_data[12]), .B1(search_data[9]), .B2(n40), 
        .C(n39), .ZN(n46) );
  AOI221D0 U15 ( .A1(n44), .A2(search_data[10]), .B1(search_data[25]), .B2(n43), .C(n42), .ZN(n45) );
  AOI221D0 U16 ( .A1(n51), .A2(search_data[7]), .B1(search_data[5]), .B2(n50), 
        .C(n49), .ZN(n65) );
  AOI221D0 U17 ( .A1(n54), .A2(search_data[16]), .B1(search_data[2]), .B2(n53), 
        .C(n52), .ZN(n64) );
  OAI221D0 U18 ( .A1(n57), .A2(search_data[3]), .B1(n56), .B2(search_data[6]), 
        .C(n55), .ZN(n62) );
  OAI221D0 U19 ( .A1(n60), .A2(search_data[1]), .B1(n59), .B2(search_data[4]), 
        .C(n58), .ZN(n61) );
  AN3D0 U20 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results)
         );
  NR2D2 U21 ( .A1(reset), .A2(n70), .ZN(n71) );
  CKND2D1 U22 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  AOI21D2 U23 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  CKND0 U24 ( .I(read_value[3]), .ZN(n57) );
  CKND0 U25 ( .I(read_value[9]), .ZN(n40) );
  CKND0 U26 ( .I(read_value[18]), .ZN(n28) );
  CKND0 U27 ( .I(read_value[6]), .ZN(n56) );
  CKND0 U28 ( .I(read_value[17]), .ZN(n24) );
  CKND0 U29 ( .I(read_value[20]), .ZN(n25) );
  CKND0 U30 ( .I(read_value[19]), .ZN(n21) );
  CKND0 U31 ( .I(read_value[22]), .ZN(n22) );
  CKND0 U32 ( .I(read_value[1]), .ZN(n60) );
  CKND0 U33 ( .I(read_value[7]), .ZN(n51) );
  CKND0 U34 ( .I(read_value[4]), .ZN(n59) );
  CKND0 U35 ( .I(read_value[16]), .ZN(n54) );
  CKND0 U36 ( .I(read_value[12]), .ZN(n41) );
  CKND0 U37 ( .I(read_value[2]), .ZN(n53) );
  CKND0 U38 ( .I(read_value[11]), .ZN(n37) );
  CKND0 U39 ( .I(read_value[14]), .ZN(n38) );
  CKND0 U40 ( .I(read_value[10]), .ZN(n44) );
  CKND0 U41 ( .I(read_value[13]), .ZN(n34) );
  CKND0 U42 ( .I(read_value[0]), .ZN(n35) );
  CKND0 U43 ( .I(read_value[25]), .ZN(n43) );
  CKND0 U44 ( .I(read_value[15]), .ZN(n27) );
  CKND0 U45 ( .I(read_value[21]), .ZN(n18) );
  CKND0 U46 ( .I(read_value[8]), .ZN(n19) );
  CKND0 U47 ( .I(read_value[23]), .ZN(n11) );
  CKND0 U48 ( .I(read_value[26]), .ZN(n12) );
  CKND0 U49 ( .I(read_value[24]), .ZN(n8) );
  CKND0 U50 ( .I(read_value[28]), .ZN(n9) );
  CKND0 U51 ( .I(read_value[27]), .ZN(n5) );
  CKND0 U52 ( .I(read_value[30]), .ZN(n6) );
  CKND0 U53 ( .I(read_value[29]), .ZN(n2) );
  CKND0 U54 ( .I(read_value[31]), .ZN(n3) );
  CKND0 U55 ( .I(read_value[5]), .ZN(n50) );
  AO22D0 U56 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U57 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U58 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U59 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U60 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U61 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U62 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U63 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U64 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U65 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U66 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U67 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U68 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U69 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U70 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U71 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U72 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U73 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U74 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U75 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  ND4D1 U76 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  NR2D1 U77 ( .A1(n62), .A2(n61), .ZN(n63) );
  AOI22D1 U78 ( .A1(search_data[1]), .A2(n60), .B1(search_data[4]), .B2(n59), 
        .ZN(n58) );
  AOI22D1 U79 ( .A1(search_data[3]), .A2(n57), .B1(search_data[6]), .B2(n56), 
        .ZN(n55) );
  OAI22D1 U80 ( .A1(n54), .A2(search_data[16]), .B1(n53), .B2(search_data[2]), 
        .ZN(n52) );
  OAI22D1 U81 ( .A1(n51), .A2(search_data[7]), .B1(n50), .B2(search_data[5]), 
        .ZN(n49) );
  ND4D1 U82 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .ZN(n67) );
  OAI22D1 U83 ( .A1(n44), .A2(search_data[10]), .B1(n43), .B2(search_data[25]), 
        .ZN(n42) );
  OAI22D1 U84 ( .A1(n41), .A2(search_data[12]), .B1(n40), .B2(search_data[9]), 
        .ZN(n39) );
  OAI22D1 U85 ( .A1(n38), .A2(search_data[14]), .B1(n37), .B2(search_data[11]), 
        .ZN(n36) );
  OAI22D1 U86 ( .A1(n35), .A2(search_data[0]), .B1(n34), .B2(search_data[13]), 
        .ZN(n33) );
  ND4D1 U87 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .ZN(n68) );
  OAI22D1 U88 ( .A1(n28), .A2(search_data[18]), .B1(n27), .B2(search_data[15]), 
        .ZN(n26) );
  OAI22D1 U89 ( .A1(n25), .A2(search_data[20]), .B1(n24), .B2(search_data[17]), 
        .ZN(n23) );
  OAI22D1 U90 ( .A1(n22), .A2(search_data[22]), .B1(n21), .B2(search_data[19]), 
        .ZN(n20) );
  OAI22D1 U91 ( .A1(n19), .A2(search_data[8]), .B1(n18), .B2(search_data[21]), 
        .ZN(n17) );
  ND4D1 U92 ( .A1(n16), .A2(n15), .A3(n14), .A4(n13), .ZN(n69) );
  OAI22D1 U93 ( .A1(n12), .A2(search_data[26]), .B1(n11), .B2(search_data[23]), 
        .ZN(n10) );
  OAI22D1 U94 ( .A1(n9), .A2(search_data[28]), .B1(n8), .B2(search_data[24]), 
        .ZN(n7) );
  OAI22D1 U95 ( .A1(n6), .A2(search_data[30]), .B1(n5), .B2(search_data[27]), 
        .ZN(n4) );
  OAI22D1 U96 ( .A1(n3), .A2(search_data[31]), .B1(n2), .B2(search_data[29]), 
        .ZN(n1) );
  AO21D1 U97 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  AO22D0 U98 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U99 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U100 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), 
        .Z(data_i[2]) );
  AO22D0 U101 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), 
        .Z(data_i[3]) );
  AO22D0 U102 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), 
        .Z(data_i[4]) );
  AO22D0 U103 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), 
        .Z(data_i[5]) );
  AO22D0 U104 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), 
        .Z(data_i[6]) );
  AO22D0 U105 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U106 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U107 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U108 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_4 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AOI221D0 U4 ( .A1(n9), .A2(search_data[31]), .B1(search_data[29]), .B2(n8), 
        .C(n7), .ZN(n22) );
  AOI221D0 U5 ( .A1(n12), .A2(search_data[30]), .B1(search_data[27]), .B2(n11), 
        .C(n10), .ZN(n21) );
  AOI221D0 U6 ( .A1(n15), .A2(search_data[28]), .B1(search_data[24]), .B2(n14), 
        .C(n13), .ZN(n20) );
  AOI221D0 U7 ( .A1(n18), .A2(search_data[26]), .B1(search_data[23]), .B2(n17), 
        .C(n16), .ZN(n19) );
  AOI221D0 U8 ( .A1(n25), .A2(search_data[8]), .B1(search_data[21]), .B2(n24), 
        .C(n23), .ZN(n38) );
  AOI221D0 U9 ( .A1(n28), .A2(search_data[22]), .B1(search_data[19]), .B2(n27), 
        .C(n26), .ZN(n37) );
  AOI221D0 U10 ( .A1(n31), .A2(search_data[20]), .B1(search_data[17]), .B2(n30), .C(n29), .ZN(n36) );
  AOI221D0 U11 ( .A1(n34), .A2(search_data[18]), .B1(search_data[15]), .B2(n33), .C(n32), .ZN(n35) );
  AOI221D0 U12 ( .A1(n41), .A2(search_data[0]), .B1(search_data[13]), .B2(n40), 
        .C(n39), .ZN(n54) );
  AOI221D0 U13 ( .A1(n44), .A2(search_data[14]), .B1(search_data[11]), .B2(n43), .C(n42), .ZN(n53) );
  AOI221D0 U14 ( .A1(n47), .A2(search_data[12]), .B1(search_data[9]), .B2(n46), 
        .C(n45), .ZN(n52) );
  AOI221D0 U15 ( .A1(n50), .A2(search_data[10]), .B1(search_data[25]), .B2(n49), .C(n48), .ZN(n51) );
  AOI221D0 U16 ( .A1(n57), .A2(search_data[7]), .B1(search_data[5]), .B2(n56), 
        .C(n55), .ZN(n65) );
  AOI221D0 U17 ( .A1(n60), .A2(search_data[16]), .B1(search_data[2]), .B2(n59), 
        .C(n58), .ZN(n64) );
  CKND0 U18 ( .I(read_value[4]), .ZN(n1) );
  CKND0 U19 ( .I(read_value[1]), .ZN(n2) );
  AOI22D0 U20 ( .A1(search_data[4]), .A2(n1), .B1(search_data[1]), .B2(n2), 
        .ZN(n3) );
  OAI221D0 U21 ( .A1(n1), .A2(search_data[4]), .B1(n2), .B2(search_data[1]), 
        .C(n3), .ZN(n61) );
  CKND0 U22 ( .I(read_value[6]), .ZN(n4) );
  CKND0 U23 ( .I(read_value[3]), .ZN(n5) );
  AOI22D0 U24 ( .A1(search_data[6]), .A2(n4), .B1(search_data[3]), .B2(n5), 
        .ZN(n6) );
  OAI221D0 U25 ( .A1(n4), .A2(search_data[6]), .B1(n5), .B2(search_data[3]), 
        .C(n6), .ZN(n62) );
  AN3D0 U26 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results)
         );
  AO21D0 U27 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U28 ( .A1(reset), .A2(n70), .ZN(n71) );
  AOI21D2 U29 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  CKND2D1 U30 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  CKND0 U31 ( .I(read_value[31]), .ZN(n9) );
  CKND0 U32 ( .I(read_value[29]), .ZN(n8) );
  CKND0 U33 ( .I(read_value[8]), .ZN(n25) );
  CKND0 U34 ( .I(read_value[21]), .ZN(n24) );
  CKND0 U35 ( .I(read_value[2]), .ZN(n59) );
  CKND0 U36 ( .I(read_value[16]), .ZN(n60) );
  CKND0 U37 ( .I(read_value[22]), .ZN(n28) );
  CKND0 U38 ( .I(read_value[5]), .ZN(n56) );
  CKND0 U39 ( .I(read_value[7]), .ZN(n57) );
  CKND0 U40 ( .I(read_value[19]), .ZN(n27) );
  CKND0 U41 ( .I(read_value[25]), .ZN(n49) );
  CKND0 U42 ( .I(read_value[10]), .ZN(n50) );
  CKND0 U43 ( .I(read_value[20]), .ZN(n31) );
  CKND0 U44 ( .I(read_value[17]), .ZN(n30) );
  CKND0 U45 ( .I(read_value[9]), .ZN(n46) );
  CKND0 U46 ( .I(read_value[12]), .ZN(n47) );
  CKND0 U47 ( .I(read_value[18]), .ZN(n34) );
  CKND0 U48 ( .I(read_value[15]), .ZN(n33) );
  CKND0 U49 ( .I(read_value[11]), .ZN(n43) );
  CKND0 U50 ( .I(read_value[14]), .ZN(n44) );
  CKND0 U51 ( .I(read_value[13]), .ZN(n40) );
  CKND0 U52 ( .I(read_value[0]), .ZN(n41) );
  CKND0 U53 ( .I(read_value[28]), .ZN(n15) );
  CKND0 U54 ( .I(read_value[24]), .ZN(n14) );
  CKND0 U55 ( .I(read_value[27]), .ZN(n11) );
  CKND0 U56 ( .I(read_value[30]), .ZN(n12) );
  CKND0 U57 ( .I(read_value[26]), .ZN(n18) );
  CKND0 U58 ( .I(read_value[23]), .ZN(n17) );
  AO22D0 U59 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), .Z(
        data_i[2]) );
  AO22D0 U60 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), .Z(
        data_i[5]) );
  AO22D0 U61 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), .Z(
        data_i[3]) );
  AO22D0 U62 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U63 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U64 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U65 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U66 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U67 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U68 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), .Z(
        data_i[4]) );
  AO22D0 U69 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U70 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U71 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U72 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), .Z(
        data_i[6]) );
  AO22D0 U73 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U74 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U75 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U76 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U77 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U78 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  ND4D1 U79 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  NR2D1 U80 ( .A1(n62), .A2(n61), .ZN(n63) );
  OAI22D1 U81 ( .A1(n60), .A2(search_data[16]), .B1(n59), .B2(search_data[2]), 
        .ZN(n58) );
  OAI22D1 U82 ( .A1(n57), .A2(search_data[7]), .B1(n56), .B2(search_data[5]), 
        .ZN(n55) );
  ND4D1 U83 ( .A1(n54), .A2(n53), .A3(n52), .A4(n51), .ZN(n67) );
  OAI22D1 U84 ( .A1(n50), .A2(search_data[10]), .B1(n49), .B2(search_data[25]), 
        .ZN(n48) );
  OAI22D1 U85 ( .A1(n47), .A2(search_data[12]), .B1(n46), .B2(search_data[9]), 
        .ZN(n45) );
  OAI22D1 U86 ( .A1(n44), .A2(search_data[14]), .B1(n43), .B2(search_data[11]), 
        .ZN(n42) );
  OAI22D1 U87 ( .A1(n41), .A2(search_data[0]), .B1(n40), .B2(search_data[13]), 
        .ZN(n39) );
  ND4D1 U88 ( .A1(n38), .A2(n37), .A3(n36), .A4(n35), .ZN(n68) );
  OAI22D1 U89 ( .A1(n34), .A2(search_data[18]), .B1(n33), .B2(search_data[15]), 
        .ZN(n32) );
  OAI22D1 U90 ( .A1(n31), .A2(search_data[20]), .B1(n30), .B2(search_data[17]), 
        .ZN(n29) );
  OAI22D1 U91 ( .A1(n28), .A2(search_data[22]), .B1(n27), .B2(search_data[19]), 
        .ZN(n26) );
  OAI22D1 U92 ( .A1(n25), .A2(search_data[8]), .B1(n24), .B2(search_data[21]), 
        .ZN(n23) );
  ND4D1 U93 ( .A1(n22), .A2(n21), .A3(n20), .A4(n19), .ZN(n69) );
  OAI22D1 U94 ( .A1(n18), .A2(search_data[26]), .B1(n17), .B2(search_data[23]), 
        .ZN(n16) );
  OAI22D1 U95 ( .A1(n15), .A2(search_data[28]), .B1(n14), .B2(search_data[24]), 
        .ZN(n13) );
  OAI22D1 U96 ( .A1(n12), .A2(search_data[30]), .B1(n11), .B2(search_data[27]), 
        .ZN(n10) );
  OAI22D1 U97 ( .A1(n9), .A2(search_data[31]), .B1(n8), .B2(search_data[29]), 
        .ZN(n7) );
  AO22D0 U98 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U99 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U100 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U101 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U102 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U103 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U104 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U105 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U106 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U107 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U108 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_5 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AOI221D0 U4 ( .A1(n9), .A2(search_data[31]), .B1(search_data[29]), .B2(n8), 
        .C(n7), .ZN(n22) );
  AOI221D0 U5 ( .A1(n12), .A2(search_data[30]), .B1(search_data[27]), .B2(n11), 
        .C(n10), .ZN(n21) );
  AOI221D0 U6 ( .A1(n15), .A2(search_data[28]), .B1(search_data[24]), .B2(n14), 
        .C(n13), .ZN(n20) );
  AOI221D0 U7 ( .A1(n18), .A2(search_data[26]), .B1(search_data[23]), .B2(n17), 
        .C(n16), .ZN(n19) );
  AOI221D0 U8 ( .A1(n25), .A2(search_data[8]), .B1(search_data[21]), .B2(n24), 
        .C(n23), .ZN(n38) );
  AOI221D0 U9 ( .A1(n28), .A2(search_data[22]), .B1(search_data[19]), .B2(n27), 
        .C(n26), .ZN(n37) );
  AOI221D0 U10 ( .A1(n31), .A2(search_data[20]), .B1(search_data[17]), .B2(n30), .C(n29), .ZN(n36) );
  AOI221D0 U11 ( .A1(n34), .A2(search_data[18]), .B1(search_data[15]), .B2(n33), .C(n32), .ZN(n35) );
  AOI221D0 U12 ( .A1(n41), .A2(search_data[0]), .B1(search_data[13]), .B2(n40), 
        .C(n39), .ZN(n54) );
  AOI221D0 U13 ( .A1(n44), .A2(search_data[14]), .B1(search_data[11]), .B2(n43), .C(n42), .ZN(n53) );
  AOI221D0 U14 ( .A1(n47), .A2(search_data[12]), .B1(search_data[9]), .B2(n46), 
        .C(n45), .ZN(n52) );
  AOI221D0 U15 ( .A1(n50), .A2(search_data[10]), .B1(search_data[25]), .B2(n49), .C(n48), .ZN(n51) );
  AOI221D0 U16 ( .A1(n57), .A2(search_data[7]), .B1(search_data[5]), .B2(n56), 
        .C(n55), .ZN(n65) );
  AOI221D0 U17 ( .A1(n60), .A2(search_data[16]), .B1(search_data[2]), .B2(n59), 
        .C(n58), .ZN(n64) );
  CKND0 U18 ( .I(read_value[4]), .ZN(n1) );
  CKND0 U19 ( .I(read_value[1]), .ZN(n2) );
  AOI22D0 U20 ( .A1(search_data[4]), .A2(n1), .B1(search_data[1]), .B2(n2), 
        .ZN(n3) );
  OAI221D0 U21 ( .A1(n1), .A2(search_data[4]), .B1(n2), .B2(search_data[1]), 
        .C(n3), .ZN(n61) );
  CKND0 U22 ( .I(read_value[6]), .ZN(n4) );
  CKND0 U23 ( .I(read_value[3]), .ZN(n5) );
  AOI22D0 U24 ( .A1(search_data[6]), .A2(n4), .B1(search_data[3]), .B2(n5), 
        .ZN(n6) );
  OAI221D0 U25 ( .A1(n4), .A2(search_data[6]), .B1(n5), .B2(search_data[3]), 
        .C(n6), .ZN(n62) );
  AN3D0 U26 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results)
         );
  AO21D0 U27 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U28 ( .A1(reset), .A2(n70), .ZN(n71) );
  CKND2D1 U29 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  AOI21D2 U30 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  CKND0 U31 ( .I(read_value[12]), .ZN(n47) );
  CKND0 U32 ( .I(read_value[9]), .ZN(n46) );
  CKND0 U33 ( .I(read_value[10]), .ZN(n50) );
  CKND0 U34 ( .I(read_value[25]), .ZN(n49) );
  CKND0 U35 ( .I(read_value[7]), .ZN(n57) );
  CKND0 U36 ( .I(read_value[5]), .ZN(n56) );
  CKND0 U37 ( .I(read_value[16]), .ZN(n60) );
  CKND0 U38 ( .I(read_value[2]), .ZN(n59) );
  CKND0 U39 ( .I(read_value[26]), .ZN(n18) );
  CKND0 U40 ( .I(read_value[23]), .ZN(n17) );
  CKND0 U41 ( .I(read_value[8]), .ZN(n25) );
  CKND0 U42 ( .I(read_value[21]), .ZN(n24) );
  CKND0 U43 ( .I(read_value[22]), .ZN(n28) );
  CKND0 U44 ( .I(read_value[19]), .ZN(n27) );
  CKND0 U45 ( .I(read_value[20]), .ZN(n31) );
  CKND0 U46 ( .I(read_value[17]), .ZN(n30) );
  CKND0 U47 ( .I(read_value[18]), .ZN(n34) );
  CKND0 U48 ( .I(read_value[15]), .ZN(n33) );
  CKND0 U49 ( .I(read_value[0]), .ZN(n41) );
  CKND0 U50 ( .I(read_value[13]), .ZN(n40) );
  CKND0 U51 ( .I(read_value[14]), .ZN(n44) );
  CKND0 U52 ( .I(read_value[11]), .ZN(n43) );
  CKND0 U53 ( .I(read_value[30]), .ZN(n12) );
  CKND0 U54 ( .I(read_value[27]), .ZN(n11) );
  CKND0 U55 ( .I(read_value[29]), .ZN(n8) );
  CKND0 U56 ( .I(read_value[31]), .ZN(n9) );
  CKND0 U57 ( .I(read_value[28]), .ZN(n15) );
  CKND0 U58 ( .I(read_value[24]), .ZN(n14) );
  AO22D0 U59 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U60 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U61 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U62 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U63 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U64 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U65 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U66 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U67 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U68 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U69 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U70 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U71 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U72 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U73 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U74 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U75 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U76 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U77 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U78 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  ND4D1 U79 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  NR2D1 U80 ( .A1(n62), .A2(n61), .ZN(n63) );
  OAI22D1 U81 ( .A1(n60), .A2(search_data[16]), .B1(n59), .B2(search_data[2]), 
        .ZN(n58) );
  OAI22D1 U82 ( .A1(n57), .A2(search_data[7]), .B1(n56), .B2(search_data[5]), 
        .ZN(n55) );
  ND4D1 U83 ( .A1(n54), .A2(n53), .A3(n52), .A4(n51), .ZN(n67) );
  OAI22D1 U84 ( .A1(n50), .A2(search_data[10]), .B1(n49), .B2(search_data[25]), 
        .ZN(n48) );
  OAI22D1 U85 ( .A1(n47), .A2(search_data[12]), .B1(n46), .B2(search_data[9]), 
        .ZN(n45) );
  OAI22D1 U86 ( .A1(n44), .A2(search_data[14]), .B1(n43), .B2(search_data[11]), 
        .ZN(n42) );
  OAI22D1 U87 ( .A1(n41), .A2(search_data[0]), .B1(n40), .B2(search_data[13]), 
        .ZN(n39) );
  ND4D1 U88 ( .A1(n38), .A2(n37), .A3(n36), .A4(n35), .ZN(n68) );
  OAI22D1 U89 ( .A1(n34), .A2(search_data[18]), .B1(n33), .B2(search_data[15]), 
        .ZN(n32) );
  OAI22D1 U90 ( .A1(n31), .A2(search_data[20]), .B1(n30), .B2(search_data[17]), 
        .ZN(n29) );
  OAI22D1 U91 ( .A1(n28), .A2(search_data[22]), .B1(n27), .B2(search_data[19]), 
        .ZN(n26) );
  OAI22D1 U92 ( .A1(n25), .A2(search_data[8]), .B1(n24), .B2(search_data[21]), 
        .ZN(n23) );
  ND4D1 U93 ( .A1(n22), .A2(n21), .A3(n20), .A4(n19), .ZN(n69) );
  OAI22D1 U94 ( .A1(n18), .A2(search_data[26]), .B1(n17), .B2(search_data[23]), 
        .ZN(n16) );
  OAI22D1 U95 ( .A1(n15), .A2(search_data[28]), .B1(n14), .B2(search_data[24]), 
        .ZN(n13) );
  OAI22D1 U96 ( .A1(n12), .A2(search_data[30]), .B1(n11), .B2(search_data[27]), 
        .ZN(n10) );
  OAI22D1 U97 ( .A1(n9), .A2(search_data[31]), .B1(n8), .B2(search_data[29]), 
        .ZN(n7) );
  AO22D0 U98 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U99 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U100 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), 
        .Z(data_i[2]) );
  AO22D0 U101 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), 
        .Z(data_i[3]) );
  AO22D0 U102 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), 
        .Z(data_i[4]) );
  AO22D0 U103 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), 
        .Z(data_i[5]) );
  AO22D0 U104 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), 
        .Z(data_i[6]) );
  AO22D0 U105 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U106 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U107 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U108 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_6 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AOI221D0 U4 ( .A1(n9), .A2(search_data[31]), .B1(search_data[29]), .B2(n8), 
        .C(n7), .ZN(n22) );
  AOI221D0 U5 ( .A1(n12), .A2(search_data[30]), .B1(search_data[27]), .B2(n11), 
        .C(n10), .ZN(n21) );
  AOI221D0 U6 ( .A1(n15), .A2(search_data[28]), .B1(search_data[24]), .B2(n14), 
        .C(n13), .ZN(n20) );
  AOI221D0 U7 ( .A1(n18), .A2(search_data[26]), .B1(search_data[23]), .B2(n17), 
        .C(n16), .ZN(n19) );
  AOI221D0 U8 ( .A1(n25), .A2(search_data[8]), .B1(search_data[21]), .B2(n24), 
        .C(n23), .ZN(n38) );
  AOI221D0 U9 ( .A1(n28), .A2(search_data[22]), .B1(search_data[19]), .B2(n27), 
        .C(n26), .ZN(n37) );
  AOI221D0 U10 ( .A1(n31), .A2(search_data[20]), .B1(search_data[17]), .B2(n30), .C(n29), .ZN(n36) );
  AOI221D0 U11 ( .A1(n34), .A2(search_data[18]), .B1(search_data[15]), .B2(n33), .C(n32), .ZN(n35) );
  AOI221D0 U12 ( .A1(n41), .A2(search_data[0]), .B1(search_data[13]), .B2(n40), 
        .C(n39), .ZN(n54) );
  AOI221D0 U13 ( .A1(n44), .A2(search_data[14]), .B1(search_data[11]), .B2(n43), .C(n42), .ZN(n53) );
  AOI221D0 U14 ( .A1(n47), .A2(search_data[12]), .B1(search_data[9]), .B2(n46), 
        .C(n45), .ZN(n52) );
  AOI221D0 U15 ( .A1(n50), .A2(search_data[10]), .B1(search_data[25]), .B2(n49), .C(n48), .ZN(n51) );
  AOI221D0 U16 ( .A1(n57), .A2(search_data[7]), .B1(search_data[5]), .B2(n56), 
        .C(n55), .ZN(n65) );
  AOI221D0 U17 ( .A1(n60), .A2(search_data[16]), .B1(search_data[2]), .B2(n59), 
        .C(n58), .ZN(n64) );
  CKND0 U18 ( .I(read_value[4]), .ZN(n1) );
  CKND0 U19 ( .I(read_value[1]), .ZN(n2) );
  AOI22D0 U20 ( .A1(search_data[4]), .A2(n1), .B1(search_data[1]), .B2(n2), 
        .ZN(n3) );
  OAI221D0 U21 ( .A1(n1), .A2(search_data[4]), .B1(n2), .B2(search_data[1]), 
        .C(n3), .ZN(n61) );
  CKND0 U22 ( .I(read_value[6]), .ZN(n4) );
  CKND0 U23 ( .I(read_value[3]), .ZN(n5) );
  AOI22D0 U24 ( .A1(search_data[6]), .A2(n4), .B1(search_data[3]), .B2(n5), 
        .ZN(n6) );
  OAI221D0 U25 ( .A1(n4), .A2(search_data[6]), .B1(n5), .B2(search_data[3]), 
        .C(n6), .ZN(n62) );
  AN3D0 U26 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results)
         );
  AO21D0 U27 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U28 ( .A1(reset), .A2(n70), .ZN(n71) );
  AOI21D2 U29 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  CKND2D1 U30 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  CKND0 U31 ( .I(read_value[30]), .ZN(n12) );
  CKND0 U32 ( .I(read_value[28]), .ZN(n15) );
  CKND0 U33 ( .I(read_value[27]), .ZN(n11) );
  CKND0 U34 ( .I(read_value[24]), .ZN(n14) );
  CKND0 U35 ( .I(read_value[26]), .ZN(n18) );
  CKND0 U36 ( .I(read_value[23]), .ZN(n17) );
  CKND0 U37 ( .I(read_value[8]), .ZN(n25) );
  CKND0 U38 ( .I(read_value[21]), .ZN(n24) );
  CKND0 U39 ( .I(read_value[31]), .ZN(n9) );
  CKND0 U40 ( .I(read_value[29]), .ZN(n8) );
  CKND0 U41 ( .I(read_value[16]), .ZN(n60) );
  CKND0 U42 ( .I(read_value[2]), .ZN(n59) );
  CKND0 U43 ( .I(read_value[22]), .ZN(n28) );
  CKND0 U44 ( .I(read_value[19]), .ZN(n27) );
  CKND0 U45 ( .I(read_value[20]), .ZN(n31) );
  CKND0 U46 ( .I(read_value[17]), .ZN(n30) );
  CKND0 U47 ( .I(read_value[18]), .ZN(n34) );
  CKND0 U48 ( .I(read_value[15]), .ZN(n33) );
  CKND0 U49 ( .I(read_value[0]), .ZN(n41) );
  CKND0 U50 ( .I(read_value[13]), .ZN(n40) );
  CKND0 U51 ( .I(read_value[14]), .ZN(n44) );
  CKND0 U52 ( .I(read_value[11]), .ZN(n43) );
  CKND0 U53 ( .I(read_value[12]), .ZN(n47) );
  CKND0 U54 ( .I(read_value[9]), .ZN(n46) );
  CKND0 U55 ( .I(read_value[10]), .ZN(n50) );
  CKND0 U56 ( .I(read_value[25]), .ZN(n49) );
  CKND0 U57 ( .I(read_value[7]), .ZN(n57) );
  CKND0 U58 ( .I(read_value[5]), .ZN(n56) );
  AO22D0 U59 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U60 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U61 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U62 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U63 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U64 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U65 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U66 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U67 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U68 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U69 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U70 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U71 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U72 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), .Z(
        data_i[6]) );
  AO22D0 U73 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), .Z(
        data_i[5]) );
  AO22D0 U74 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), .Z(
        data_i[4]) );
  AO22D0 U75 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), .Z(
        data_i[3]) );
  AO22D0 U76 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), .Z(
        data_i[2]) );
  AO22D0 U77 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U78 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  ND4D1 U79 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  NR2D1 U80 ( .A1(n62), .A2(n61), .ZN(n63) );
  OAI22D1 U81 ( .A1(n60), .A2(search_data[16]), .B1(n59), .B2(search_data[2]), 
        .ZN(n58) );
  OAI22D1 U82 ( .A1(n57), .A2(search_data[7]), .B1(n56), .B2(search_data[5]), 
        .ZN(n55) );
  ND4D1 U83 ( .A1(n54), .A2(n53), .A3(n52), .A4(n51), .ZN(n67) );
  OAI22D1 U84 ( .A1(n50), .A2(search_data[10]), .B1(n49), .B2(search_data[25]), 
        .ZN(n48) );
  OAI22D1 U85 ( .A1(n47), .A2(search_data[12]), .B1(n46), .B2(search_data[9]), 
        .ZN(n45) );
  OAI22D1 U86 ( .A1(n44), .A2(search_data[14]), .B1(n43), .B2(search_data[11]), 
        .ZN(n42) );
  OAI22D1 U87 ( .A1(n41), .A2(search_data[0]), .B1(n40), .B2(search_data[13]), 
        .ZN(n39) );
  ND4D1 U88 ( .A1(n38), .A2(n37), .A3(n36), .A4(n35), .ZN(n68) );
  OAI22D1 U89 ( .A1(n34), .A2(search_data[18]), .B1(n33), .B2(search_data[15]), 
        .ZN(n32) );
  OAI22D1 U90 ( .A1(n31), .A2(search_data[20]), .B1(n30), .B2(search_data[17]), 
        .ZN(n29) );
  OAI22D1 U91 ( .A1(n28), .A2(search_data[22]), .B1(n27), .B2(search_data[19]), 
        .ZN(n26) );
  OAI22D1 U92 ( .A1(n25), .A2(search_data[8]), .B1(n24), .B2(search_data[21]), 
        .ZN(n23) );
  ND4D1 U93 ( .A1(n22), .A2(n21), .A3(n20), .A4(n19), .ZN(n69) );
  OAI22D1 U94 ( .A1(n18), .A2(search_data[26]), .B1(n17), .B2(search_data[23]), 
        .ZN(n16) );
  OAI22D1 U95 ( .A1(n15), .A2(search_data[28]), .B1(n14), .B2(search_data[24]), 
        .ZN(n13) );
  OAI22D1 U96 ( .A1(n12), .A2(search_data[30]), .B1(n11), .B2(search_data[27]), 
        .ZN(n10) );
  OAI22D1 U97 ( .A1(n9), .A2(search_data[31]), .B1(n8), .B2(search_data[29]), 
        .ZN(n7) );
  AO22D0 U98 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U99 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U100 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U101 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U102 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U103 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U104 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U105 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U106 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U107 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U108 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_7 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AOI221D0 U4 ( .A1(n3), .A2(search_data[31]), .B1(search_data[29]), .B2(n2), 
        .C(n1), .ZN(n16) );
  AOI221D0 U5 ( .A1(n6), .A2(search_data[30]), .B1(search_data[27]), .B2(n5), 
        .C(n4), .ZN(n15) );
  AOI221D0 U6 ( .A1(n9), .A2(search_data[28]), .B1(search_data[24]), .B2(n8), 
        .C(n7), .ZN(n14) );
  AOI221D0 U7 ( .A1(n12), .A2(search_data[26]), .B1(search_data[23]), .B2(n11), 
        .C(n10), .ZN(n13) );
  AOI221D0 U8 ( .A1(n19), .A2(search_data[8]), .B1(search_data[21]), .B2(n18), 
        .C(n17), .ZN(n32) );
  AOI221D0 U9 ( .A1(n22), .A2(search_data[22]), .B1(search_data[19]), .B2(n21), 
        .C(n20), .ZN(n31) );
  AOI221D0 U10 ( .A1(n25), .A2(search_data[20]), .B1(search_data[17]), .B2(n24), .C(n23), .ZN(n30) );
  AOI221D0 U11 ( .A1(n28), .A2(search_data[18]), .B1(search_data[15]), .B2(n27), .C(n26), .ZN(n29) );
  AOI221D0 U12 ( .A1(n35), .A2(search_data[0]), .B1(search_data[13]), .B2(n34), 
        .C(n33), .ZN(n48) );
  AOI221D0 U13 ( .A1(n38), .A2(search_data[14]), .B1(search_data[11]), .B2(n37), .C(n36), .ZN(n47) );
  AOI221D0 U14 ( .A1(n41), .A2(search_data[12]), .B1(search_data[9]), .B2(n40), 
        .C(n39), .ZN(n46) );
  AOI221D0 U15 ( .A1(n44), .A2(search_data[10]), .B1(search_data[25]), .B2(n43), .C(n42), .ZN(n45) );
  AOI221D0 U16 ( .A1(n51), .A2(search_data[7]), .B1(search_data[5]), .B2(n50), 
        .C(n49), .ZN(n65) );
  AOI221D0 U17 ( .A1(n54), .A2(search_data[16]), .B1(search_data[2]), .B2(n53), 
        .C(n52), .ZN(n64) );
  OAI221D0 U18 ( .A1(n57), .A2(search_data[3]), .B1(n56), .B2(search_data[6]), 
        .C(n55), .ZN(n62) );
  OAI221D0 U19 ( .A1(n60), .A2(search_data[1]), .B1(n59), .B2(search_data[4]), 
        .C(n58), .ZN(n61) );
  AN3D0 U20 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results)
         );
  AO21D0 U21 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U22 ( .A1(reset), .A2(n70), .ZN(n71) );
  AOI21D2 U23 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  CKND2D1 U24 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  CKND0 U25 ( .I(read_value[2]), .ZN(n53) );
  CKND0 U26 ( .I(read_value[16]), .ZN(n54) );
  CKND0 U27 ( .I(read_value[5]), .ZN(n50) );
  CKND0 U28 ( .I(read_value[7]), .ZN(n51) );
  CKND0 U29 ( .I(read_value[4]), .ZN(n59) );
  CKND0 U30 ( .I(read_value[1]), .ZN(n60) );
  CKND0 U31 ( .I(read_value[6]), .ZN(n56) );
  CKND0 U32 ( .I(read_value[3]), .ZN(n57) );
  CKND0 U33 ( .I(read_value[13]), .ZN(n34) );
  CKND0 U34 ( .I(read_value[0]), .ZN(n35) );
  CKND0 U35 ( .I(read_value[15]), .ZN(n27) );
  CKND0 U36 ( .I(read_value[18]), .ZN(n28) );
  CKND0 U37 ( .I(read_value[31]), .ZN(n3) );
  CKND0 U38 ( .I(read_value[29]), .ZN(n2) );
  CKND0 U39 ( .I(read_value[30]), .ZN(n6) );
  CKND0 U40 ( .I(read_value[17]), .ZN(n24) );
  CKND0 U41 ( .I(read_value[27]), .ZN(n5) );
  CKND0 U42 ( .I(read_value[20]), .ZN(n25) );
  CKND0 U43 ( .I(read_value[28]), .ZN(n9) );
  CKND0 U44 ( .I(read_value[24]), .ZN(n8) );
  CKND0 U45 ( .I(read_value[26]), .ZN(n12) );
  CKND0 U46 ( .I(read_value[23]), .ZN(n11) );
  CKND0 U47 ( .I(read_value[19]), .ZN(n21) );
  CKND0 U48 ( .I(read_value[22]), .ZN(n22) );
  CKND0 U49 ( .I(read_value[8]), .ZN(n19) );
  CKND0 U50 ( .I(read_value[21]), .ZN(n18) );
  CKND0 U51 ( .I(read_value[25]), .ZN(n43) );
  CKND0 U52 ( .I(read_value[10]), .ZN(n44) );
  CKND0 U53 ( .I(read_value[9]), .ZN(n40) );
  CKND0 U54 ( .I(read_value[12]), .ZN(n41) );
  CKND0 U55 ( .I(read_value[11]), .ZN(n37) );
  CKND0 U56 ( .I(read_value[14]), .ZN(n38) );
  AO22D0 U57 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U58 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U59 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U60 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U61 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U62 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U63 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U64 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U65 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U66 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U67 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U68 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U69 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U70 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U71 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U72 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U73 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U74 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U75 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U76 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  ND4D1 U77 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  NR2D1 U78 ( .A1(n62), .A2(n61), .ZN(n63) );
  AOI22D1 U79 ( .A1(search_data[1]), .A2(n60), .B1(search_data[4]), .B2(n59), 
        .ZN(n58) );
  AOI22D1 U80 ( .A1(search_data[3]), .A2(n57), .B1(search_data[6]), .B2(n56), 
        .ZN(n55) );
  OAI22D1 U81 ( .A1(n54), .A2(search_data[16]), .B1(n53), .B2(search_data[2]), 
        .ZN(n52) );
  OAI22D1 U82 ( .A1(n51), .A2(search_data[7]), .B1(n50), .B2(search_data[5]), 
        .ZN(n49) );
  ND4D1 U83 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .ZN(n67) );
  OAI22D1 U84 ( .A1(n44), .A2(search_data[10]), .B1(n43), .B2(search_data[25]), 
        .ZN(n42) );
  OAI22D1 U85 ( .A1(n41), .A2(search_data[12]), .B1(n40), .B2(search_data[9]), 
        .ZN(n39) );
  OAI22D1 U86 ( .A1(n38), .A2(search_data[14]), .B1(n37), .B2(search_data[11]), 
        .ZN(n36) );
  OAI22D1 U87 ( .A1(n35), .A2(search_data[0]), .B1(n34), .B2(search_data[13]), 
        .ZN(n33) );
  ND4D1 U88 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .ZN(n68) );
  OAI22D1 U89 ( .A1(n28), .A2(search_data[18]), .B1(n27), .B2(search_data[15]), 
        .ZN(n26) );
  OAI22D1 U90 ( .A1(n25), .A2(search_data[20]), .B1(n24), .B2(search_data[17]), 
        .ZN(n23) );
  OAI22D1 U91 ( .A1(n22), .A2(search_data[22]), .B1(n21), .B2(search_data[19]), 
        .ZN(n20) );
  OAI22D1 U92 ( .A1(n19), .A2(search_data[8]), .B1(n18), .B2(search_data[21]), 
        .ZN(n17) );
  ND4D1 U93 ( .A1(n16), .A2(n15), .A3(n14), .A4(n13), .ZN(n69) );
  OAI22D1 U94 ( .A1(n12), .A2(search_data[26]), .B1(n11), .B2(search_data[23]), 
        .ZN(n10) );
  OAI22D1 U95 ( .A1(n9), .A2(search_data[28]), .B1(n8), .B2(search_data[24]), 
        .ZN(n7) );
  OAI22D1 U96 ( .A1(n6), .A2(search_data[30]), .B1(n5), .B2(search_data[27]), 
        .ZN(n4) );
  OAI22D1 U97 ( .A1(n3), .A2(search_data[31]), .B1(n2), .B2(search_data[29]), 
        .ZN(n1) );
  AO22D0 U98 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U99 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U100 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), 
        .Z(data_i[2]) );
  AO22D0 U101 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), 
        .Z(data_i[3]) );
  AO22D0 U102 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), 
        .Z(data_i[4]) );
  AO22D0 U103 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), 
        .Z(data_i[5]) );
  AO22D0 U104 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), 
        .Z(data_i[6]) );
  AO22D0 U105 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U106 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U107 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U108 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_8 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AOI221D0 U4 ( .A1(n9), .A2(search_data[31]), .B1(search_data[29]), .B2(n8), 
        .C(n7), .ZN(n22) );
  AOI221D0 U5 ( .A1(n12), .A2(search_data[30]), .B1(search_data[27]), .B2(n11), 
        .C(n10), .ZN(n21) );
  AOI221D0 U6 ( .A1(n15), .A2(search_data[28]), .B1(search_data[24]), .B2(n14), 
        .C(n13), .ZN(n20) );
  AOI221D0 U7 ( .A1(n18), .A2(search_data[26]), .B1(search_data[23]), .B2(n17), 
        .C(n16), .ZN(n19) );
  AOI221D0 U8 ( .A1(n25), .A2(search_data[8]), .B1(search_data[21]), .B2(n24), 
        .C(n23), .ZN(n38) );
  AOI221D0 U9 ( .A1(n28), .A2(search_data[22]), .B1(search_data[19]), .B2(n27), 
        .C(n26), .ZN(n37) );
  AOI221D0 U10 ( .A1(n31), .A2(search_data[20]), .B1(search_data[17]), .B2(n30), .C(n29), .ZN(n36) );
  AOI221D0 U11 ( .A1(n34), .A2(search_data[18]), .B1(search_data[15]), .B2(n33), .C(n32), .ZN(n35) );
  AOI221D0 U12 ( .A1(n41), .A2(search_data[0]), .B1(search_data[13]), .B2(n40), 
        .C(n39), .ZN(n54) );
  AOI221D0 U13 ( .A1(n44), .A2(search_data[14]), .B1(search_data[11]), .B2(n43), .C(n42), .ZN(n53) );
  AOI221D0 U14 ( .A1(n47), .A2(search_data[12]), .B1(search_data[9]), .B2(n46), 
        .C(n45), .ZN(n52) );
  AOI221D0 U15 ( .A1(n50), .A2(search_data[10]), .B1(search_data[25]), .B2(n49), .C(n48), .ZN(n51) );
  AOI221D0 U16 ( .A1(n57), .A2(search_data[7]), .B1(search_data[5]), .B2(n56), 
        .C(n55), .ZN(n65) );
  AOI221D0 U17 ( .A1(n60), .A2(search_data[16]), .B1(search_data[2]), .B2(n59), 
        .C(n58), .ZN(n64) );
  CKND0 U18 ( .I(read_value[4]), .ZN(n1) );
  CKND0 U19 ( .I(read_value[1]), .ZN(n2) );
  AOI22D0 U20 ( .A1(search_data[4]), .A2(n1), .B1(search_data[1]), .B2(n2), 
        .ZN(n3) );
  OAI221D0 U21 ( .A1(n1), .A2(search_data[4]), .B1(n2), .B2(search_data[1]), 
        .C(n3), .ZN(n61) );
  CKND0 U22 ( .I(read_value[6]), .ZN(n4) );
  CKND0 U23 ( .I(read_value[3]), .ZN(n5) );
  AOI22D0 U24 ( .A1(search_data[6]), .A2(n4), .B1(search_data[3]), .B2(n5), 
        .ZN(n6) );
  OAI221D0 U25 ( .A1(n4), .A2(search_data[6]), .B1(n5), .B2(search_data[3]), 
        .C(n6), .ZN(n62) );
  AN3D0 U26 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results)
         );
  AO21D0 U27 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U28 ( .A1(reset), .A2(n70), .ZN(n71) );
  CKND2D1 U29 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  AOI21D2 U30 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  CKND0 U31 ( .I(read_value[2]), .ZN(n59) );
  CKND0 U32 ( .I(read_value[16]), .ZN(n60) );
  CKND0 U33 ( .I(read_value[5]), .ZN(n56) );
  CKND0 U34 ( .I(read_value[7]), .ZN(n57) );
  CKND0 U35 ( .I(read_value[19]), .ZN(n27) );
  CKND0 U36 ( .I(read_value[22]), .ZN(n28) );
  CKND0 U37 ( .I(read_value[21]), .ZN(n24) );
  CKND0 U38 ( .I(read_value[8]), .ZN(n25) );
  CKND0 U39 ( .I(read_value[23]), .ZN(n17) );
  CKND0 U40 ( .I(read_value[26]), .ZN(n18) );
  CKND0 U41 ( .I(read_value[24]), .ZN(n14) );
  CKND0 U42 ( .I(read_value[28]), .ZN(n15) );
  CKND0 U43 ( .I(read_value[27]), .ZN(n11) );
  CKND0 U44 ( .I(read_value[30]), .ZN(n12) );
  CKND0 U45 ( .I(read_value[29]), .ZN(n8) );
  CKND0 U46 ( .I(read_value[31]), .ZN(n9) );
  CKND0 U47 ( .I(read_value[25]), .ZN(n49) );
  CKND0 U48 ( .I(read_value[10]), .ZN(n50) );
  CKND0 U49 ( .I(read_value[9]), .ZN(n46) );
  CKND0 U50 ( .I(read_value[12]), .ZN(n47) );
  CKND0 U51 ( .I(read_value[11]), .ZN(n43) );
  CKND0 U52 ( .I(read_value[14]), .ZN(n44) );
  CKND0 U53 ( .I(read_value[13]), .ZN(n40) );
  CKND0 U54 ( .I(read_value[0]), .ZN(n41) );
  CKND0 U55 ( .I(read_value[15]), .ZN(n33) );
  CKND0 U56 ( .I(read_value[18]), .ZN(n34) );
  CKND0 U57 ( .I(read_value[17]), .ZN(n30) );
  CKND0 U58 ( .I(read_value[20]), .ZN(n31) );
  AO22D0 U59 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U60 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U61 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U62 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U63 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U64 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U65 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U66 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U67 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U68 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U69 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U70 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U71 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U72 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U73 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U74 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U75 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U76 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U77 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U78 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  ND4D1 U79 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  NR2D1 U80 ( .A1(n62), .A2(n61), .ZN(n63) );
  OAI22D1 U81 ( .A1(n60), .A2(search_data[16]), .B1(n59), .B2(search_data[2]), 
        .ZN(n58) );
  OAI22D1 U82 ( .A1(n57), .A2(search_data[7]), .B1(n56), .B2(search_data[5]), 
        .ZN(n55) );
  ND4D1 U83 ( .A1(n54), .A2(n53), .A3(n52), .A4(n51), .ZN(n67) );
  OAI22D1 U84 ( .A1(n50), .A2(search_data[10]), .B1(n49), .B2(search_data[25]), 
        .ZN(n48) );
  OAI22D1 U85 ( .A1(n47), .A2(search_data[12]), .B1(n46), .B2(search_data[9]), 
        .ZN(n45) );
  OAI22D1 U86 ( .A1(n44), .A2(search_data[14]), .B1(n43), .B2(search_data[11]), 
        .ZN(n42) );
  OAI22D1 U87 ( .A1(n41), .A2(search_data[0]), .B1(n40), .B2(search_data[13]), 
        .ZN(n39) );
  ND4D1 U88 ( .A1(n38), .A2(n37), .A3(n36), .A4(n35), .ZN(n68) );
  OAI22D1 U89 ( .A1(n34), .A2(search_data[18]), .B1(n33), .B2(search_data[15]), 
        .ZN(n32) );
  OAI22D1 U90 ( .A1(n31), .A2(search_data[20]), .B1(n30), .B2(search_data[17]), 
        .ZN(n29) );
  OAI22D1 U91 ( .A1(n28), .A2(search_data[22]), .B1(n27), .B2(search_data[19]), 
        .ZN(n26) );
  OAI22D1 U92 ( .A1(n25), .A2(search_data[8]), .B1(n24), .B2(search_data[21]), 
        .ZN(n23) );
  ND4D1 U93 ( .A1(n22), .A2(n21), .A3(n20), .A4(n19), .ZN(n69) );
  OAI22D1 U94 ( .A1(n18), .A2(search_data[26]), .B1(n17), .B2(search_data[23]), 
        .ZN(n16) );
  OAI22D1 U95 ( .A1(n15), .A2(search_data[28]), .B1(n14), .B2(search_data[24]), 
        .ZN(n13) );
  OAI22D1 U96 ( .A1(n12), .A2(search_data[30]), .B1(n11), .B2(search_data[27]), 
        .ZN(n10) );
  OAI22D1 U97 ( .A1(n9), .A2(search_data[31]), .B1(n8), .B2(search_data[29]), 
        .ZN(n7) );
  AO22D0 U98 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U99 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U100 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), 
        .Z(data_i[2]) );
  AO22D0 U101 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), 
        .Z(data_i[3]) );
  AO22D0 U102 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), 
        .Z(data_i[4]) );
  AO22D0 U103 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), 
        .Z(data_i[5]) );
  AO22D0 U104 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), 
        .Z(data_i[6]) );
  AO22D0 U105 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U106 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U107 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U108 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_9 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AOI221D0 U4 ( .A1(n9), .A2(search_data[31]), .B1(search_data[29]), .B2(n8), 
        .C(n7), .ZN(n22) );
  AOI221D0 U5 ( .A1(n12), .A2(search_data[30]), .B1(search_data[27]), .B2(n11), 
        .C(n10), .ZN(n21) );
  AOI221D0 U6 ( .A1(n15), .A2(search_data[28]), .B1(search_data[24]), .B2(n14), 
        .C(n13), .ZN(n20) );
  AOI221D0 U7 ( .A1(n18), .A2(search_data[26]), .B1(search_data[23]), .B2(n17), 
        .C(n16), .ZN(n19) );
  AOI221D0 U8 ( .A1(n25), .A2(search_data[8]), .B1(search_data[21]), .B2(n24), 
        .C(n23), .ZN(n38) );
  AOI221D0 U9 ( .A1(n28), .A2(search_data[22]), .B1(search_data[19]), .B2(n27), 
        .C(n26), .ZN(n37) );
  AOI221D0 U10 ( .A1(n31), .A2(search_data[20]), .B1(search_data[17]), .B2(n30), .C(n29), .ZN(n36) );
  AOI221D0 U11 ( .A1(n34), .A2(search_data[18]), .B1(search_data[15]), .B2(n33), .C(n32), .ZN(n35) );
  AOI221D0 U12 ( .A1(n41), .A2(search_data[0]), .B1(search_data[13]), .B2(n40), 
        .C(n39), .ZN(n54) );
  AOI221D0 U13 ( .A1(n44), .A2(search_data[14]), .B1(search_data[11]), .B2(n43), .C(n42), .ZN(n53) );
  AOI221D0 U14 ( .A1(n47), .A2(search_data[12]), .B1(search_data[9]), .B2(n46), 
        .C(n45), .ZN(n52) );
  AOI221D0 U15 ( .A1(n50), .A2(search_data[10]), .B1(search_data[25]), .B2(n49), .C(n48), .ZN(n51) );
  AOI221D0 U16 ( .A1(n57), .A2(search_data[7]), .B1(search_data[5]), .B2(n56), 
        .C(n55), .ZN(n65) );
  AOI221D0 U17 ( .A1(n60), .A2(search_data[16]), .B1(search_data[2]), .B2(n59), 
        .C(n58), .ZN(n64) );
  CKND0 U18 ( .I(read_value[4]), .ZN(n1) );
  CKND0 U19 ( .I(read_value[1]), .ZN(n2) );
  AOI22D0 U20 ( .A1(search_data[4]), .A2(n1), .B1(search_data[1]), .B2(n2), 
        .ZN(n3) );
  OAI221D0 U21 ( .A1(n1), .A2(search_data[4]), .B1(n2), .B2(search_data[1]), 
        .C(n3), .ZN(n61) );
  CKND0 U22 ( .I(read_value[6]), .ZN(n4) );
  CKND0 U23 ( .I(read_value[3]), .ZN(n5) );
  AOI22D0 U24 ( .A1(search_data[6]), .A2(n4), .B1(search_data[3]), .B2(n5), 
        .ZN(n6) );
  OAI221D0 U25 ( .A1(n4), .A2(search_data[6]), .B1(n5), .B2(search_data[3]), 
        .C(n6), .ZN(n62) );
  AN3D0 U26 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results)
         );
  AO21D0 U27 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U28 ( .A1(reset), .A2(n70), .ZN(n71) );
  AOI21D2 U29 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  CKND2D1 U30 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  CKND0 U31 ( .I(read_value[31]), .ZN(n9) );
  CKND0 U32 ( .I(read_value[0]), .ZN(n41) );
  CKND0 U33 ( .I(read_value[13]), .ZN(n40) );
  CKND0 U34 ( .I(read_value[14]), .ZN(n44) );
  CKND0 U35 ( .I(read_value[11]), .ZN(n43) );
  CKND0 U36 ( .I(read_value[12]), .ZN(n47) );
  CKND0 U37 ( .I(read_value[9]), .ZN(n46) );
  CKND0 U38 ( .I(read_value[10]), .ZN(n50) );
  CKND0 U39 ( .I(read_value[25]), .ZN(n49) );
  CKND0 U40 ( .I(read_value[7]), .ZN(n57) );
  CKND0 U41 ( .I(read_value[5]), .ZN(n56) );
  CKND0 U42 ( .I(read_value[16]), .ZN(n60) );
  CKND0 U43 ( .I(read_value[2]), .ZN(n59) );
  CKND0 U44 ( .I(read_value[29]), .ZN(n8) );
  CKND0 U45 ( .I(read_value[30]), .ZN(n12) );
  CKND0 U46 ( .I(read_value[27]), .ZN(n11) );
  CKND0 U47 ( .I(read_value[28]), .ZN(n15) );
  CKND0 U48 ( .I(read_value[24]), .ZN(n14) );
  CKND0 U49 ( .I(read_value[26]), .ZN(n18) );
  CKND0 U50 ( .I(read_value[23]), .ZN(n17) );
  CKND0 U51 ( .I(read_value[8]), .ZN(n25) );
  CKND0 U52 ( .I(read_value[21]), .ZN(n24) );
  CKND0 U53 ( .I(read_value[22]), .ZN(n28) );
  CKND0 U54 ( .I(read_value[19]), .ZN(n27) );
  CKND0 U55 ( .I(read_value[20]), .ZN(n31) );
  CKND0 U56 ( .I(read_value[17]), .ZN(n30) );
  CKND0 U57 ( .I(read_value[18]), .ZN(n34) );
  CKND0 U58 ( .I(read_value[15]), .ZN(n33) );
  AO22D0 U59 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U60 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U61 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U62 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U63 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U64 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U65 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U66 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U67 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), .Z(
        data_i[6]) );
  AO22D0 U68 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U69 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U70 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U71 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), .Z(
        data_i[5]) );
  AO22D0 U72 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U73 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U74 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), .Z(
        data_i[3]) );
  AO22D0 U75 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), .Z(
        data_i[2]) );
  AO22D0 U76 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U77 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U78 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), .Z(
        data_i[4]) );
  ND4D1 U79 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  NR2D1 U80 ( .A1(n62), .A2(n61), .ZN(n63) );
  OAI22D1 U81 ( .A1(n60), .A2(search_data[16]), .B1(n59), .B2(search_data[2]), 
        .ZN(n58) );
  OAI22D1 U82 ( .A1(n57), .A2(search_data[7]), .B1(n56), .B2(search_data[5]), 
        .ZN(n55) );
  ND4D1 U83 ( .A1(n54), .A2(n53), .A3(n52), .A4(n51), .ZN(n67) );
  OAI22D1 U84 ( .A1(n50), .A2(search_data[10]), .B1(n49), .B2(search_data[25]), 
        .ZN(n48) );
  OAI22D1 U85 ( .A1(n47), .A2(search_data[12]), .B1(n46), .B2(search_data[9]), 
        .ZN(n45) );
  OAI22D1 U86 ( .A1(n44), .A2(search_data[14]), .B1(n43), .B2(search_data[11]), 
        .ZN(n42) );
  OAI22D1 U87 ( .A1(n41), .A2(search_data[0]), .B1(n40), .B2(search_data[13]), 
        .ZN(n39) );
  ND4D1 U88 ( .A1(n38), .A2(n37), .A3(n36), .A4(n35), .ZN(n68) );
  OAI22D1 U89 ( .A1(n34), .A2(search_data[18]), .B1(n33), .B2(search_data[15]), 
        .ZN(n32) );
  OAI22D1 U90 ( .A1(n31), .A2(search_data[20]), .B1(n30), .B2(search_data[17]), 
        .ZN(n29) );
  OAI22D1 U91 ( .A1(n28), .A2(search_data[22]), .B1(n27), .B2(search_data[19]), 
        .ZN(n26) );
  OAI22D1 U92 ( .A1(n25), .A2(search_data[8]), .B1(n24), .B2(search_data[21]), 
        .ZN(n23) );
  ND4D1 U93 ( .A1(n22), .A2(n21), .A3(n20), .A4(n19), .ZN(n69) );
  OAI22D1 U94 ( .A1(n18), .A2(search_data[26]), .B1(n17), .B2(search_data[23]), 
        .ZN(n16) );
  OAI22D1 U95 ( .A1(n15), .A2(search_data[28]), .B1(n14), .B2(search_data[24]), 
        .ZN(n13) );
  OAI22D1 U96 ( .A1(n12), .A2(search_data[30]), .B1(n11), .B2(search_data[27]), 
        .ZN(n10) );
  OAI22D1 U97 ( .A1(n9), .A2(search_data[31]), .B1(n8), .B2(search_data[29]), 
        .ZN(n7) );
  AO22D0 U98 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U99 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U100 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U101 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U102 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U103 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U104 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U105 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U106 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U107 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U108 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_10 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AOI221D0 U4 ( .A1(n3), .A2(search_data[31]), .B1(search_data[29]), .B2(n2), 
        .C(n1), .ZN(n16) );
  AOI221D0 U5 ( .A1(n6), .A2(search_data[30]), .B1(search_data[27]), .B2(n5), 
        .C(n4), .ZN(n15) );
  AOI221D0 U6 ( .A1(n9), .A2(search_data[28]), .B1(search_data[24]), .B2(n8), 
        .C(n7), .ZN(n14) );
  AOI221D0 U7 ( .A1(n12), .A2(search_data[26]), .B1(search_data[23]), .B2(n11), 
        .C(n10), .ZN(n13) );
  AOI221D0 U8 ( .A1(n19), .A2(search_data[8]), .B1(search_data[21]), .B2(n18), 
        .C(n17), .ZN(n32) );
  AOI221D0 U9 ( .A1(n22), .A2(search_data[22]), .B1(search_data[19]), .B2(n21), 
        .C(n20), .ZN(n31) );
  AOI221D0 U10 ( .A1(n25), .A2(search_data[20]), .B1(search_data[17]), .B2(n24), .C(n23), .ZN(n30) );
  AOI221D0 U11 ( .A1(n28), .A2(search_data[18]), .B1(search_data[15]), .B2(n27), .C(n26), .ZN(n29) );
  AOI221D0 U12 ( .A1(n35), .A2(search_data[0]), .B1(search_data[13]), .B2(n34), 
        .C(n33), .ZN(n48) );
  AOI221D0 U13 ( .A1(n38), .A2(search_data[14]), .B1(search_data[11]), .B2(n37), .C(n36), .ZN(n47) );
  AOI221D0 U14 ( .A1(n41), .A2(search_data[12]), .B1(search_data[9]), .B2(n40), 
        .C(n39), .ZN(n46) );
  AOI221D0 U15 ( .A1(n44), .A2(search_data[10]), .B1(search_data[25]), .B2(n43), .C(n42), .ZN(n45) );
  AOI221D0 U16 ( .A1(n51), .A2(search_data[7]), .B1(search_data[5]), .B2(n50), 
        .C(n49), .ZN(n65) );
  AOI221D0 U17 ( .A1(n54), .A2(search_data[16]), .B1(search_data[2]), .B2(n53), 
        .C(n52), .ZN(n64) );
  OAI221D0 U18 ( .A1(n57), .A2(search_data[3]), .B1(n56), .B2(search_data[6]), 
        .C(n55), .ZN(n62) );
  OAI221D0 U19 ( .A1(n60), .A2(search_data[1]), .B1(n59), .B2(search_data[4]), 
        .C(n58), .ZN(n61) );
  AN3D0 U20 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results)
         );
  AO21D0 U21 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U22 ( .A1(reset), .A2(n70), .ZN(n71) );
  AOI21D2 U23 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  CKND2D1 U24 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  CKND0 U25 ( .I(read_value[26]), .ZN(n12) );
  CKND0 U26 ( .I(read_value[5]), .ZN(n50) );
  CKND0 U27 ( .I(read_value[23]), .ZN(n11) );
  CKND0 U28 ( .I(read_value[7]), .ZN(n51) );
  CKND0 U29 ( .I(read_value[8]), .ZN(n19) );
  CKND0 U30 ( .I(read_value[25]), .ZN(n43) );
  CKND0 U31 ( .I(read_value[21]), .ZN(n18) );
  CKND0 U32 ( .I(read_value[10]), .ZN(n44) );
  CKND0 U33 ( .I(read_value[22]), .ZN(n22) );
  CKND0 U34 ( .I(read_value[9]), .ZN(n40) );
  CKND0 U35 ( .I(read_value[12]), .ZN(n41) );
  CKND0 U36 ( .I(read_value[19]), .ZN(n21) );
  CKND0 U37 ( .I(read_value[11]), .ZN(n37) );
  CKND0 U38 ( .I(read_value[20]), .ZN(n25) );
  CKND0 U39 ( .I(read_value[14]), .ZN(n38) );
  CKND0 U40 ( .I(read_value[17]), .ZN(n24) );
  CKND0 U41 ( .I(read_value[13]), .ZN(n34) );
  CKND0 U42 ( .I(read_value[18]), .ZN(n28) );
  CKND0 U43 ( .I(read_value[0]), .ZN(n35) );
  CKND0 U44 ( .I(read_value[15]), .ZN(n27) );
  CKND0 U45 ( .I(read_value[31]), .ZN(n3) );
  CKND0 U46 ( .I(read_value[29]), .ZN(n2) );
  CKND0 U47 ( .I(read_value[4]), .ZN(n59) );
  CKND0 U48 ( .I(read_value[1]), .ZN(n60) );
  CKND0 U49 ( .I(read_value[30]), .ZN(n6) );
  CKND0 U50 ( .I(read_value[27]), .ZN(n5) );
  CKND0 U51 ( .I(read_value[6]), .ZN(n56) );
  CKND0 U52 ( .I(read_value[3]), .ZN(n57) );
  CKND0 U53 ( .I(read_value[28]), .ZN(n9) );
  CKND0 U54 ( .I(read_value[2]), .ZN(n53) );
  CKND0 U55 ( .I(read_value[24]), .ZN(n8) );
  CKND0 U56 ( .I(read_value[16]), .ZN(n54) );
  AO22D0 U57 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U58 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U59 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U60 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U61 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U62 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U63 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U64 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U65 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U66 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U67 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U68 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U69 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U70 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), .Z(
        data_i[6]) );
  AO22D0 U71 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), .Z(
        data_i[5]) );
  AO22D0 U72 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), .Z(
        data_i[4]) );
  AO22D0 U73 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), .Z(
        data_i[3]) );
  AO22D0 U74 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), .Z(
        data_i[2]) );
  AO22D0 U75 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U76 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  ND4D1 U77 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  NR2D1 U78 ( .A1(n62), .A2(n61), .ZN(n63) );
  AOI22D1 U79 ( .A1(search_data[1]), .A2(n60), .B1(search_data[4]), .B2(n59), 
        .ZN(n58) );
  AOI22D1 U80 ( .A1(search_data[3]), .A2(n57), .B1(search_data[6]), .B2(n56), 
        .ZN(n55) );
  OAI22D1 U81 ( .A1(n54), .A2(search_data[16]), .B1(n53), .B2(search_data[2]), 
        .ZN(n52) );
  OAI22D1 U82 ( .A1(n51), .A2(search_data[7]), .B1(n50), .B2(search_data[5]), 
        .ZN(n49) );
  ND4D1 U83 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .ZN(n67) );
  OAI22D1 U84 ( .A1(n44), .A2(search_data[10]), .B1(n43), .B2(search_data[25]), 
        .ZN(n42) );
  OAI22D1 U85 ( .A1(n41), .A2(search_data[12]), .B1(n40), .B2(search_data[9]), 
        .ZN(n39) );
  OAI22D1 U86 ( .A1(n38), .A2(search_data[14]), .B1(n37), .B2(search_data[11]), 
        .ZN(n36) );
  OAI22D1 U87 ( .A1(n35), .A2(search_data[0]), .B1(n34), .B2(search_data[13]), 
        .ZN(n33) );
  ND4D1 U88 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .ZN(n68) );
  OAI22D1 U89 ( .A1(n28), .A2(search_data[18]), .B1(n27), .B2(search_data[15]), 
        .ZN(n26) );
  OAI22D1 U90 ( .A1(n25), .A2(search_data[20]), .B1(n24), .B2(search_data[17]), 
        .ZN(n23) );
  OAI22D1 U91 ( .A1(n22), .A2(search_data[22]), .B1(n21), .B2(search_data[19]), 
        .ZN(n20) );
  OAI22D1 U92 ( .A1(n19), .A2(search_data[8]), .B1(n18), .B2(search_data[21]), 
        .ZN(n17) );
  ND4D1 U93 ( .A1(n16), .A2(n15), .A3(n14), .A4(n13), .ZN(n69) );
  OAI22D1 U94 ( .A1(n12), .A2(search_data[26]), .B1(n11), .B2(search_data[23]), 
        .ZN(n10) );
  OAI22D1 U95 ( .A1(n9), .A2(search_data[28]), .B1(n8), .B2(search_data[24]), 
        .ZN(n7) );
  OAI22D1 U96 ( .A1(n6), .A2(search_data[30]), .B1(n5), .B2(search_data[27]), 
        .ZN(n4) );
  OAI22D1 U97 ( .A1(n3), .A2(search_data[31]), .B1(n2), .B2(search_data[29]), 
        .ZN(n1) );
  AO22D0 U98 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U99 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U100 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U101 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U102 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U103 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U104 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U105 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U106 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U107 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U108 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_11 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AOI221D0 U4 ( .A1(n3), .A2(search_data[31]), .B1(search_data[29]), .B2(n2), 
        .C(n1), .ZN(n16) );
  AOI221D0 U5 ( .A1(n6), .A2(search_data[30]), .B1(search_data[27]), .B2(n5), 
        .C(n4), .ZN(n15) );
  AOI221D0 U6 ( .A1(n9), .A2(search_data[28]), .B1(search_data[24]), .B2(n8), 
        .C(n7), .ZN(n14) );
  AOI221D0 U7 ( .A1(n12), .A2(search_data[26]), .B1(search_data[23]), .B2(n11), 
        .C(n10), .ZN(n13) );
  AOI221D0 U8 ( .A1(n19), .A2(search_data[8]), .B1(search_data[21]), .B2(n18), 
        .C(n17), .ZN(n32) );
  AOI221D0 U9 ( .A1(n22), .A2(search_data[22]), .B1(search_data[19]), .B2(n21), 
        .C(n20), .ZN(n31) );
  AOI221D0 U10 ( .A1(n25), .A2(search_data[20]), .B1(search_data[17]), .B2(n24), .C(n23), .ZN(n30) );
  AOI221D0 U11 ( .A1(n28), .A2(search_data[18]), .B1(search_data[15]), .B2(n27), .C(n26), .ZN(n29) );
  AOI221D0 U12 ( .A1(n35), .A2(search_data[0]), .B1(search_data[13]), .B2(n34), 
        .C(n33), .ZN(n48) );
  AOI221D0 U13 ( .A1(n38), .A2(search_data[14]), .B1(search_data[11]), .B2(n37), .C(n36), .ZN(n47) );
  AOI221D0 U14 ( .A1(n41), .A2(search_data[12]), .B1(search_data[9]), .B2(n40), 
        .C(n39), .ZN(n46) );
  AOI221D0 U15 ( .A1(n44), .A2(search_data[10]), .B1(search_data[25]), .B2(n43), .C(n42), .ZN(n45) );
  AOI221D0 U16 ( .A1(n51), .A2(search_data[7]), .B1(search_data[5]), .B2(n50), 
        .C(n49), .ZN(n65) );
  AOI221D0 U17 ( .A1(n54), .A2(search_data[16]), .B1(search_data[2]), .B2(n53), 
        .C(n52), .ZN(n64) );
  OAI221D0 U18 ( .A1(n57), .A2(search_data[3]), .B1(n56), .B2(search_data[6]), 
        .C(n55), .ZN(n62) );
  OAI221D0 U19 ( .A1(n60), .A2(search_data[1]), .B1(n59), .B2(search_data[4]), 
        .C(n58), .ZN(n61) );
  AN3D0 U20 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results)
         );
  AO21D0 U21 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U22 ( .A1(reset), .A2(n70), .ZN(n71) );
  CKND2D1 U23 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  AOI21D2 U24 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  CKND0 U25 ( .I(read_value[15]), .ZN(n27) );
  CKND0 U26 ( .I(read_value[18]), .ZN(n28) );
  CKND0 U27 ( .I(read_value[17]), .ZN(n24) );
  CKND0 U28 ( .I(read_value[20]), .ZN(n25) );
  CKND0 U29 ( .I(read_value[19]), .ZN(n21) );
  CKND0 U30 ( .I(read_value[22]), .ZN(n22) );
  CKND0 U31 ( .I(read_value[21]), .ZN(n18) );
  CKND0 U32 ( .I(read_value[8]), .ZN(n19) );
  CKND0 U33 ( .I(read_value[23]), .ZN(n11) );
  CKND0 U34 ( .I(read_value[26]), .ZN(n12) );
  CKND0 U35 ( .I(read_value[24]), .ZN(n8) );
  CKND0 U36 ( .I(read_value[7]), .ZN(n51) );
  CKND0 U37 ( .I(read_value[25]), .ZN(n43) );
  CKND0 U38 ( .I(read_value[10]), .ZN(n44) );
  CKND0 U39 ( .I(read_value[9]), .ZN(n40) );
  CKND0 U40 ( .I(read_value[12]), .ZN(n41) );
  CKND0 U41 ( .I(read_value[5]), .ZN(n50) );
  CKND0 U42 ( .I(read_value[11]), .ZN(n37) );
  CKND0 U43 ( .I(read_value[14]), .ZN(n38) );
  CKND0 U44 ( .I(read_value[13]), .ZN(n34) );
  CKND0 U45 ( .I(read_value[0]), .ZN(n35) );
  CKND0 U46 ( .I(read_value[28]), .ZN(n9) );
  CKND0 U47 ( .I(read_value[27]), .ZN(n5) );
  CKND0 U48 ( .I(read_value[30]), .ZN(n6) );
  CKND0 U49 ( .I(read_value[29]), .ZN(n2) );
  CKND0 U50 ( .I(read_value[31]), .ZN(n3) );
  CKND0 U51 ( .I(read_value[4]), .ZN(n59) );
  CKND0 U52 ( .I(read_value[2]), .ZN(n53) );
  CKND0 U53 ( .I(read_value[16]), .ZN(n54) );
  CKND0 U54 ( .I(read_value[3]), .ZN(n57) );
  CKND0 U55 ( .I(read_value[1]), .ZN(n60) );
  CKND0 U56 ( .I(read_value[6]), .ZN(n56) );
  AO22D0 U57 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U58 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U59 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U60 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), .Z(
        data_i[2]) );
  AO22D0 U61 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), .Z(
        data_i[3]) );
  AO22D0 U62 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), .Z(
        data_i[4]) );
  AO22D0 U63 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), .Z(
        data_i[5]) );
  AO22D0 U64 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), .Z(
        data_i[6]) );
  AO22D0 U65 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U66 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U67 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U68 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U69 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U70 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U71 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U72 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U73 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U74 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U75 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U76 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  ND4D1 U77 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  NR2D1 U78 ( .A1(n62), .A2(n61), .ZN(n63) );
  AOI22D1 U79 ( .A1(search_data[1]), .A2(n60), .B1(search_data[4]), .B2(n59), 
        .ZN(n58) );
  AOI22D1 U80 ( .A1(search_data[3]), .A2(n57), .B1(search_data[6]), .B2(n56), 
        .ZN(n55) );
  OAI22D1 U81 ( .A1(n54), .A2(search_data[16]), .B1(n53), .B2(search_data[2]), 
        .ZN(n52) );
  OAI22D1 U82 ( .A1(n51), .A2(search_data[7]), .B1(n50), .B2(search_data[5]), 
        .ZN(n49) );
  ND4D1 U83 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .ZN(n67) );
  OAI22D1 U84 ( .A1(n44), .A2(search_data[10]), .B1(n43), .B2(search_data[25]), 
        .ZN(n42) );
  OAI22D1 U85 ( .A1(n41), .A2(search_data[12]), .B1(n40), .B2(search_data[9]), 
        .ZN(n39) );
  OAI22D1 U86 ( .A1(n38), .A2(search_data[14]), .B1(n37), .B2(search_data[11]), 
        .ZN(n36) );
  OAI22D1 U87 ( .A1(n35), .A2(search_data[0]), .B1(n34), .B2(search_data[13]), 
        .ZN(n33) );
  ND4D1 U88 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .ZN(n68) );
  OAI22D1 U89 ( .A1(n28), .A2(search_data[18]), .B1(n27), .B2(search_data[15]), 
        .ZN(n26) );
  OAI22D1 U90 ( .A1(n25), .A2(search_data[20]), .B1(n24), .B2(search_data[17]), 
        .ZN(n23) );
  OAI22D1 U91 ( .A1(n22), .A2(search_data[22]), .B1(n21), .B2(search_data[19]), 
        .ZN(n20) );
  OAI22D1 U92 ( .A1(n19), .A2(search_data[8]), .B1(n18), .B2(search_data[21]), 
        .ZN(n17) );
  ND4D1 U93 ( .A1(n16), .A2(n15), .A3(n14), .A4(n13), .ZN(n69) );
  OAI22D1 U94 ( .A1(n12), .A2(search_data[26]), .B1(n11), .B2(search_data[23]), 
        .ZN(n10) );
  OAI22D1 U95 ( .A1(n9), .A2(search_data[28]), .B1(n8), .B2(search_data[24]), 
        .ZN(n7) );
  OAI22D1 U96 ( .A1(n6), .A2(search_data[30]), .B1(n5), .B2(search_data[27]), 
        .ZN(n4) );
  OAI22D1 U97 ( .A1(n3), .A2(search_data[31]), .B1(n2), .B2(search_data[29]), 
        .ZN(n1) );
  AO22D0 U98 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U99 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U100 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U101 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U102 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U103 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U104 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U105 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U106 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U107 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U108 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_12 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AOI221D0 U4 ( .A1(n9), .A2(search_data[31]), .B1(search_data[29]), .B2(n8), 
        .C(n7), .ZN(n22) );
  AOI221D0 U5 ( .A1(n12), .A2(search_data[30]), .B1(search_data[27]), .B2(n11), 
        .C(n10), .ZN(n21) );
  AOI221D0 U6 ( .A1(n15), .A2(search_data[28]), .B1(search_data[24]), .B2(n14), 
        .C(n13), .ZN(n20) );
  AOI221D0 U7 ( .A1(n18), .A2(search_data[26]), .B1(search_data[23]), .B2(n17), 
        .C(n16), .ZN(n19) );
  AOI221D0 U8 ( .A1(n25), .A2(search_data[8]), .B1(search_data[21]), .B2(n24), 
        .C(n23), .ZN(n38) );
  AOI221D0 U9 ( .A1(n28), .A2(search_data[22]), .B1(search_data[19]), .B2(n27), 
        .C(n26), .ZN(n37) );
  AOI221D0 U10 ( .A1(n31), .A2(search_data[20]), .B1(search_data[17]), .B2(n30), .C(n29), .ZN(n36) );
  AOI221D0 U11 ( .A1(n34), .A2(search_data[18]), .B1(search_data[15]), .B2(n33), .C(n32), .ZN(n35) );
  AOI221D0 U12 ( .A1(n41), .A2(search_data[0]), .B1(search_data[13]), .B2(n40), 
        .C(n39), .ZN(n54) );
  AOI221D0 U13 ( .A1(n44), .A2(search_data[14]), .B1(search_data[11]), .B2(n43), .C(n42), .ZN(n53) );
  AOI221D0 U14 ( .A1(n47), .A2(search_data[12]), .B1(search_data[9]), .B2(n46), 
        .C(n45), .ZN(n52) );
  AOI221D0 U15 ( .A1(n50), .A2(search_data[10]), .B1(search_data[25]), .B2(n49), .C(n48), .ZN(n51) );
  AOI221D0 U16 ( .A1(n57), .A2(search_data[7]), .B1(search_data[5]), .B2(n56), 
        .C(n55), .ZN(n65) );
  AOI221D0 U17 ( .A1(n60), .A2(search_data[16]), .B1(search_data[2]), .B2(n59), 
        .C(n58), .ZN(n64) );
  CKND0 U18 ( .I(read_value[4]), .ZN(n1) );
  CKND0 U19 ( .I(read_value[1]), .ZN(n2) );
  AOI22D0 U20 ( .A1(search_data[4]), .A2(n1), .B1(search_data[1]), .B2(n2), 
        .ZN(n3) );
  OAI221D0 U21 ( .A1(n1), .A2(search_data[4]), .B1(n2), .B2(search_data[1]), 
        .C(n3), .ZN(n61) );
  CKND0 U22 ( .I(read_value[6]), .ZN(n4) );
  CKND0 U23 ( .I(read_value[3]), .ZN(n5) );
  AOI22D0 U24 ( .A1(search_data[6]), .A2(n4), .B1(search_data[3]), .B2(n5), 
        .ZN(n6) );
  OAI221D0 U25 ( .A1(n4), .A2(search_data[6]), .B1(n5), .B2(search_data[3]), 
        .C(n6), .ZN(n62) );
  AN3D0 U26 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results)
         );
  AO21D0 U27 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U28 ( .A1(reset), .A2(n70), .ZN(n71) );
  AOI21D2 U29 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  CKND2D1 U30 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  CKND0 U31 ( .I(read_value[13]), .ZN(n40) );
  CKND0 U32 ( .I(read_value[16]), .ZN(n60) );
  CKND0 U33 ( .I(read_value[9]), .ZN(n46) );
  CKND0 U34 ( .I(read_value[2]), .ZN(n59) );
  CKND0 U35 ( .I(read_value[0]), .ZN(n41) );
  CKND0 U36 ( .I(read_value[25]), .ZN(n49) );
  CKND0 U37 ( .I(read_value[10]), .ZN(n50) );
  CKND0 U38 ( .I(read_value[11]), .ZN(n43) );
  CKND0 U39 ( .I(read_value[12]), .ZN(n47) );
  CKND0 U40 ( .I(read_value[14]), .ZN(n44) );
  CKND0 U41 ( .I(read_value[7]), .ZN(n57) );
  CKND0 U42 ( .I(read_value[5]), .ZN(n56) );
  CKND0 U43 ( .I(read_value[28]), .ZN(n15) );
  CKND0 U44 ( .I(read_value[24]), .ZN(n14) );
  CKND0 U45 ( .I(read_value[17]), .ZN(n30) );
  CKND0 U46 ( .I(read_value[26]), .ZN(n18) );
  CKND0 U47 ( .I(read_value[23]), .ZN(n17) );
  CKND0 U48 ( .I(read_value[20]), .ZN(n31) );
  CKND0 U49 ( .I(read_value[8]), .ZN(n25) );
  CKND0 U50 ( .I(read_value[21]), .ZN(n24) );
  CKND0 U51 ( .I(read_value[19]), .ZN(n27) );
  CKND0 U52 ( .I(read_value[22]), .ZN(n28) );
  CKND0 U53 ( .I(read_value[31]), .ZN(n9) );
  CKND0 U54 ( .I(read_value[29]), .ZN(n8) );
  CKND0 U55 ( .I(read_value[15]), .ZN(n33) );
  CKND0 U56 ( .I(read_value[30]), .ZN(n12) );
  CKND0 U57 ( .I(read_value[18]), .ZN(n34) );
  CKND0 U58 ( .I(read_value[27]), .ZN(n11) );
  AO22D0 U59 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U60 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U61 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U62 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U63 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U64 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U65 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U66 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U67 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U68 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U69 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U70 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U71 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U72 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U73 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U74 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U75 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U76 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U77 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U78 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  ND4D1 U79 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  NR2D1 U80 ( .A1(n62), .A2(n61), .ZN(n63) );
  OAI22D1 U81 ( .A1(n60), .A2(search_data[16]), .B1(n59), .B2(search_data[2]), 
        .ZN(n58) );
  OAI22D1 U82 ( .A1(n57), .A2(search_data[7]), .B1(n56), .B2(search_data[5]), 
        .ZN(n55) );
  ND4D1 U83 ( .A1(n54), .A2(n53), .A3(n52), .A4(n51), .ZN(n67) );
  OAI22D1 U84 ( .A1(n50), .A2(search_data[10]), .B1(n49), .B2(search_data[25]), 
        .ZN(n48) );
  OAI22D1 U85 ( .A1(n47), .A2(search_data[12]), .B1(n46), .B2(search_data[9]), 
        .ZN(n45) );
  OAI22D1 U86 ( .A1(n44), .A2(search_data[14]), .B1(n43), .B2(search_data[11]), 
        .ZN(n42) );
  OAI22D1 U87 ( .A1(n41), .A2(search_data[0]), .B1(n40), .B2(search_data[13]), 
        .ZN(n39) );
  ND4D1 U88 ( .A1(n38), .A2(n37), .A3(n36), .A4(n35), .ZN(n68) );
  OAI22D1 U89 ( .A1(n34), .A2(search_data[18]), .B1(n33), .B2(search_data[15]), 
        .ZN(n32) );
  OAI22D1 U90 ( .A1(n31), .A2(search_data[20]), .B1(n30), .B2(search_data[17]), 
        .ZN(n29) );
  OAI22D1 U91 ( .A1(n28), .A2(search_data[22]), .B1(n27), .B2(search_data[19]), 
        .ZN(n26) );
  OAI22D1 U92 ( .A1(n25), .A2(search_data[8]), .B1(n24), .B2(search_data[21]), 
        .ZN(n23) );
  ND4D1 U93 ( .A1(n22), .A2(n21), .A3(n20), .A4(n19), .ZN(n69) );
  OAI22D1 U94 ( .A1(n18), .A2(search_data[26]), .B1(n17), .B2(search_data[23]), 
        .ZN(n16) );
  OAI22D1 U95 ( .A1(n15), .A2(search_data[28]), .B1(n14), .B2(search_data[24]), 
        .ZN(n13) );
  OAI22D1 U96 ( .A1(n12), .A2(search_data[30]), .B1(n11), .B2(search_data[27]), 
        .ZN(n10) );
  OAI22D1 U97 ( .A1(n9), .A2(search_data[31]), .B1(n8), .B2(search_data[29]), 
        .ZN(n7) );
  AO22D0 U98 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U99 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U100 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), 
        .Z(data_i[2]) );
  AO22D0 U101 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), 
        .Z(data_i[3]) );
  AO22D0 U102 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), 
        .Z(data_i[4]) );
  AO22D0 U103 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), 
        .Z(data_i[5]) );
  AO22D0 U104 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), 
        .Z(data_i[6]) );
  AO22D0 U105 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U106 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U107 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U108 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_13 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AOI221D0 U4 ( .A1(n9), .A2(search_data[31]), .B1(search_data[29]), .B2(n8), 
        .C(n7), .ZN(n22) );
  AOI221D0 U5 ( .A1(n12), .A2(search_data[30]), .B1(search_data[27]), .B2(n11), 
        .C(n10), .ZN(n21) );
  AOI221D0 U6 ( .A1(n15), .A2(search_data[28]), .B1(search_data[24]), .B2(n14), 
        .C(n13), .ZN(n20) );
  AOI221D0 U7 ( .A1(n18), .A2(search_data[26]), .B1(search_data[23]), .B2(n17), 
        .C(n16), .ZN(n19) );
  AOI221D0 U8 ( .A1(n25), .A2(search_data[8]), .B1(search_data[21]), .B2(n24), 
        .C(n23), .ZN(n38) );
  AOI221D0 U9 ( .A1(n28), .A2(search_data[22]), .B1(search_data[19]), .B2(n27), 
        .C(n26), .ZN(n37) );
  AOI221D0 U10 ( .A1(n31), .A2(search_data[20]), .B1(search_data[17]), .B2(n30), .C(n29), .ZN(n36) );
  AOI221D0 U11 ( .A1(n34), .A2(search_data[18]), .B1(search_data[15]), .B2(n33), .C(n32), .ZN(n35) );
  AOI221D0 U12 ( .A1(n41), .A2(search_data[0]), .B1(search_data[13]), .B2(n40), 
        .C(n39), .ZN(n54) );
  AOI221D0 U13 ( .A1(n44), .A2(search_data[14]), .B1(search_data[11]), .B2(n43), .C(n42), .ZN(n53) );
  AOI221D0 U14 ( .A1(n47), .A2(search_data[12]), .B1(search_data[9]), .B2(n46), 
        .C(n45), .ZN(n52) );
  AOI221D0 U15 ( .A1(n50), .A2(search_data[10]), .B1(search_data[25]), .B2(n49), .C(n48), .ZN(n51) );
  AOI221D0 U16 ( .A1(n57), .A2(search_data[7]), .B1(search_data[5]), .B2(n56), 
        .C(n55), .ZN(n65) );
  AOI221D0 U17 ( .A1(n60), .A2(search_data[16]), .B1(search_data[2]), .B2(n59), 
        .C(n58), .ZN(n64) );
  CKND0 U18 ( .I(read_value[4]), .ZN(n1) );
  CKND0 U19 ( .I(read_value[1]), .ZN(n2) );
  AOI22D0 U20 ( .A1(search_data[4]), .A2(n1), .B1(search_data[1]), .B2(n2), 
        .ZN(n3) );
  OAI221D0 U21 ( .A1(n1), .A2(search_data[4]), .B1(n2), .B2(search_data[1]), 
        .C(n3), .ZN(n61) );
  CKND0 U22 ( .I(read_value[6]), .ZN(n4) );
  CKND0 U23 ( .I(read_value[3]), .ZN(n5) );
  AOI22D0 U24 ( .A1(search_data[6]), .A2(n4), .B1(search_data[3]), .B2(n5), 
        .ZN(n6) );
  OAI221D0 U25 ( .A1(n4), .A2(search_data[6]), .B1(n5), .B2(search_data[3]), 
        .C(n6), .ZN(n62) );
  AN3D0 U26 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results)
         );
  AO21D0 U27 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U28 ( .A1(reset), .A2(n70), .ZN(n71) );
  AOI21D2 U29 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  CKND2D1 U30 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  CKND0 U31 ( .I(read_value[7]), .ZN(n57) );
  CKND0 U32 ( .I(read_value[5]), .ZN(n56) );
  CKND0 U33 ( .I(read_value[25]), .ZN(n49) );
  CKND0 U34 ( .I(read_value[10]), .ZN(n50) );
  CKND0 U35 ( .I(read_value[9]), .ZN(n46) );
  CKND0 U36 ( .I(read_value[2]), .ZN(n59) );
  CKND0 U37 ( .I(read_value[16]), .ZN(n60) );
  CKND0 U38 ( .I(read_value[19]), .ZN(n27) );
  CKND0 U39 ( .I(read_value[22]), .ZN(n28) );
  CKND0 U40 ( .I(read_value[31]), .ZN(n9) );
  CKND0 U41 ( .I(read_value[21]), .ZN(n24) );
  CKND0 U42 ( .I(read_value[8]), .ZN(n25) );
  CKND0 U43 ( .I(read_value[29]), .ZN(n8) );
  CKND0 U44 ( .I(read_value[23]), .ZN(n17) );
  CKND0 U45 ( .I(read_value[26]), .ZN(n18) );
  CKND0 U46 ( .I(read_value[24]), .ZN(n14) );
  CKND0 U47 ( .I(read_value[30]), .ZN(n12) );
  CKND0 U48 ( .I(read_value[28]), .ZN(n15) );
  CKND0 U49 ( .I(read_value[27]), .ZN(n11) );
  CKND0 U50 ( .I(read_value[12]), .ZN(n47) );
  CKND0 U51 ( .I(read_value[11]), .ZN(n43) );
  CKND0 U52 ( .I(read_value[14]), .ZN(n44) );
  CKND0 U53 ( .I(read_value[13]), .ZN(n40) );
  CKND0 U54 ( .I(read_value[0]), .ZN(n41) );
  CKND0 U55 ( .I(read_value[15]), .ZN(n33) );
  CKND0 U56 ( .I(read_value[18]), .ZN(n34) );
  CKND0 U57 ( .I(read_value[17]), .ZN(n30) );
  CKND0 U58 ( .I(read_value[20]), .ZN(n31) );
  AO22D0 U59 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U60 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U61 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U62 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U63 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U64 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U65 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U66 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U67 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U68 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U69 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U70 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U71 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U72 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U73 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U74 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U75 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U76 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U77 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U78 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  ND4D1 U79 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  NR2D1 U80 ( .A1(n62), .A2(n61), .ZN(n63) );
  OAI22D1 U81 ( .A1(n60), .A2(search_data[16]), .B1(n59), .B2(search_data[2]), 
        .ZN(n58) );
  OAI22D1 U82 ( .A1(n57), .A2(search_data[7]), .B1(n56), .B2(search_data[5]), 
        .ZN(n55) );
  ND4D1 U83 ( .A1(n54), .A2(n53), .A3(n52), .A4(n51), .ZN(n67) );
  OAI22D1 U84 ( .A1(n50), .A2(search_data[10]), .B1(n49), .B2(search_data[25]), 
        .ZN(n48) );
  OAI22D1 U85 ( .A1(n47), .A2(search_data[12]), .B1(n46), .B2(search_data[9]), 
        .ZN(n45) );
  OAI22D1 U86 ( .A1(n44), .A2(search_data[14]), .B1(n43), .B2(search_data[11]), 
        .ZN(n42) );
  OAI22D1 U87 ( .A1(n41), .A2(search_data[0]), .B1(n40), .B2(search_data[13]), 
        .ZN(n39) );
  ND4D1 U88 ( .A1(n38), .A2(n37), .A3(n36), .A4(n35), .ZN(n68) );
  OAI22D1 U89 ( .A1(n34), .A2(search_data[18]), .B1(n33), .B2(search_data[15]), 
        .ZN(n32) );
  OAI22D1 U90 ( .A1(n31), .A2(search_data[20]), .B1(n30), .B2(search_data[17]), 
        .ZN(n29) );
  OAI22D1 U91 ( .A1(n28), .A2(search_data[22]), .B1(n27), .B2(search_data[19]), 
        .ZN(n26) );
  OAI22D1 U92 ( .A1(n25), .A2(search_data[8]), .B1(n24), .B2(search_data[21]), 
        .ZN(n23) );
  ND4D1 U93 ( .A1(n22), .A2(n21), .A3(n20), .A4(n19), .ZN(n69) );
  OAI22D1 U94 ( .A1(n18), .A2(search_data[26]), .B1(n17), .B2(search_data[23]), 
        .ZN(n16) );
  OAI22D1 U95 ( .A1(n15), .A2(search_data[28]), .B1(n14), .B2(search_data[24]), 
        .ZN(n13) );
  OAI22D1 U96 ( .A1(n12), .A2(search_data[30]), .B1(n11), .B2(search_data[27]), 
        .ZN(n10) );
  OAI22D1 U97 ( .A1(n9), .A2(search_data[31]), .B1(n8), .B2(search_data[29]), 
        .ZN(n7) );
  AO22D0 U98 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U99 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U100 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), 
        .Z(data_i[2]) );
  AO22D0 U101 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), 
        .Z(data_i[3]) );
  AO22D0 U102 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), 
        .Z(data_i[4]) );
  AO22D0 U103 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), 
        .Z(data_i[5]) );
  AO22D0 U104 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), 
        .Z(data_i[6]) );
  AO22D0 U105 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U106 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U107 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U108 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_14 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AOI221D0 U4 ( .A1(n3), .A2(search_data[31]), .B1(search_data[29]), .B2(n2), 
        .C(n1), .ZN(n16) );
  AOI221D0 U5 ( .A1(n6), .A2(search_data[30]), .B1(search_data[27]), .B2(n5), 
        .C(n4), .ZN(n15) );
  AOI221D0 U6 ( .A1(n9), .A2(search_data[28]), .B1(search_data[24]), .B2(n8), 
        .C(n7), .ZN(n14) );
  AOI221D0 U7 ( .A1(n12), .A2(search_data[26]), .B1(search_data[23]), .B2(n11), 
        .C(n10), .ZN(n13) );
  AOI221D0 U8 ( .A1(n19), .A2(search_data[8]), .B1(search_data[21]), .B2(n18), 
        .C(n17), .ZN(n32) );
  AOI221D0 U9 ( .A1(n22), .A2(search_data[22]), .B1(search_data[19]), .B2(n21), 
        .C(n20), .ZN(n31) );
  AOI221D0 U10 ( .A1(n25), .A2(search_data[20]), .B1(search_data[17]), .B2(n24), .C(n23), .ZN(n30) );
  AOI221D0 U11 ( .A1(n28), .A2(search_data[18]), .B1(search_data[15]), .B2(n27), .C(n26), .ZN(n29) );
  AOI221D0 U12 ( .A1(n35), .A2(search_data[0]), .B1(search_data[13]), .B2(n34), 
        .C(n33), .ZN(n48) );
  AOI221D0 U13 ( .A1(n38), .A2(search_data[14]), .B1(search_data[11]), .B2(n37), .C(n36), .ZN(n47) );
  AOI221D0 U14 ( .A1(n41), .A2(search_data[12]), .B1(search_data[9]), .B2(n40), 
        .C(n39), .ZN(n46) );
  AOI221D0 U15 ( .A1(n44), .A2(search_data[10]), .B1(search_data[25]), .B2(n43), .C(n42), .ZN(n45) );
  AOI221D0 U16 ( .A1(n51), .A2(search_data[7]), .B1(search_data[5]), .B2(n50), 
        .C(n49), .ZN(n65) );
  AOI221D0 U17 ( .A1(n54), .A2(search_data[16]), .B1(search_data[2]), .B2(n53), 
        .C(n52), .ZN(n64) );
  OAI221D0 U18 ( .A1(n57), .A2(search_data[3]), .B1(n56), .B2(search_data[6]), 
        .C(n55), .ZN(n62) );
  OAI221D0 U19 ( .A1(n60), .A2(search_data[1]), .B1(n59), .B2(search_data[4]), 
        .C(n58), .ZN(n61) );
  AN3D0 U20 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results)
         );
  AO21D0 U21 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U22 ( .A1(reset), .A2(n70), .ZN(n71) );
  AOI21D2 U23 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  CKND2D1 U24 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  CKND0 U25 ( .I(read_value[17]), .ZN(n24) );
  CKND0 U26 ( .I(read_value[15]), .ZN(n27) );
  CKND0 U27 ( .I(read_value[18]), .ZN(n28) );
  CKND0 U28 ( .I(read_value[9]), .ZN(n40) );
  CKND0 U29 ( .I(read_value[11]), .ZN(n37) );
  CKND0 U30 ( .I(read_value[14]), .ZN(n38) );
  CKND0 U31 ( .I(read_value[12]), .ZN(n41) );
  CKND0 U32 ( .I(read_value[13]), .ZN(n34) );
  CKND0 U33 ( .I(read_value[0]), .ZN(n35) );
  CKND0 U34 ( .I(read_value[23]), .ZN(n11) );
  CKND0 U35 ( .I(read_value[31]), .ZN(n3) );
  CKND0 U36 ( .I(read_value[26]), .ZN(n12) );
  CKND0 U37 ( .I(read_value[29]), .ZN(n2) );
  CKND0 U38 ( .I(read_value[24]), .ZN(n8) );
  CKND0 U39 ( .I(read_value[28]), .ZN(n9) );
  CKND0 U40 ( .I(read_value[27]), .ZN(n5) );
  CKND0 U41 ( .I(read_value[30]), .ZN(n6) );
  CKND0 U42 ( .I(read_value[20]), .ZN(n25) );
  CKND0 U43 ( .I(read_value[19]), .ZN(n21) );
  CKND0 U44 ( .I(read_value[22]), .ZN(n22) );
  CKND0 U45 ( .I(read_value[21]), .ZN(n18) );
  CKND0 U46 ( .I(read_value[8]), .ZN(n19) );
  CKND0 U47 ( .I(read_value[5]), .ZN(n50) );
  CKND0 U48 ( .I(read_value[16]), .ZN(n54) );
  CKND0 U49 ( .I(read_value[2]), .ZN(n53) );
  CKND0 U50 ( .I(read_value[3]), .ZN(n57) );
  CKND0 U51 ( .I(read_value[6]), .ZN(n56) );
  CKND0 U52 ( .I(read_value[4]), .ZN(n59) );
  CKND0 U53 ( .I(read_value[1]), .ZN(n60) );
  CKND0 U54 ( .I(read_value[25]), .ZN(n43) );
  CKND0 U55 ( .I(read_value[10]), .ZN(n44) );
  CKND0 U56 ( .I(read_value[7]), .ZN(n51) );
  AO22D0 U57 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U58 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U59 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U60 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U61 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U62 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U63 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U64 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U65 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U66 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U67 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U68 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U69 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U70 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U71 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U72 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U73 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U74 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U75 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U76 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  ND4D1 U77 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  NR2D1 U78 ( .A1(n62), .A2(n61), .ZN(n63) );
  AOI22D1 U79 ( .A1(search_data[1]), .A2(n60), .B1(search_data[4]), .B2(n59), 
        .ZN(n58) );
  AOI22D1 U80 ( .A1(search_data[3]), .A2(n57), .B1(search_data[6]), .B2(n56), 
        .ZN(n55) );
  OAI22D1 U81 ( .A1(n54), .A2(search_data[16]), .B1(n53), .B2(search_data[2]), 
        .ZN(n52) );
  OAI22D1 U82 ( .A1(n51), .A2(search_data[7]), .B1(n50), .B2(search_data[5]), 
        .ZN(n49) );
  ND4D1 U83 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .ZN(n67) );
  OAI22D1 U84 ( .A1(n44), .A2(search_data[10]), .B1(n43), .B2(search_data[25]), 
        .ZN(n42) );
  OAI22D1 U85 ( .A1(n41), .A2(search_data[12]), .B1(n40), .B2(search_data[9]), 
        .ZN(n39) );
  OAI22D1 U86 ( .A1(n38), .A2(search_data[14]), .B1(n37), .B2(search_data[11]), 
        .ZN(n36) );
  OAI22D1 U87 ( .A1(n35), .A2(search_data[0]), .B1(n34), .B2(search_data[13]), 
        .ZN(n33) );
  ND4D1 U88 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .ZN(n68) );
  OAI22D1 U89 ( .A1(n28), .A2(search_data[18]), .B1(n27), .B2(search_data[15]), 
        .ZN(n26) );
  OAI22D1 U90 ( .A1(n25), .A2(search_data[20]), .B1(n24), .B2(search_data[17]), 
        .ZN(n23) );
  OAI22D1 U91 ( .A1(n22), .A2(search_data[22]), .B1(n21), .B2(search_data[19]), 
        .ZN(n20) );
  OAI22D1 U92 ( .A1(n19), .A2(search_data[8]), .B1(n18), .B2(search_data[21]), 
        .ZN(n17) );
  ND4D1 U93 ( .A1(n16), .A2(n15), .A3(n14), .A4(n13), .ZN(n69) );
  OAI22D1 U94 ( .A1(n12), .A2(search_data[26]), .B1(n11), .B2(search_data[23]), 
        .ZN(n10) );
  OAI22D1 U95 ( .A1(n9), .A2(search_data[28]), .B1(n8), .B2(search_data[24]), 
        .ZN(n7) );
  OAI22D1 U96 ( .A1(n6), .A2(search_data[30]), .B1(n5), .B2(search_data[27]), 
        .ZN(n4) );
  OAI22D1 U97 ( .A1(n3), .A2(search_data[31]), .B1(n2), .B2(search_data[29]), 
        .ZN(n1) );
  AO22D0 U98 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U99 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U100 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), 
        .Z(data_i[2]) );
  AO22D0 U101 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), 
        .Z(data_i[3]) );
  AO22D0 U102 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), 
        .Z(data_i[4]) );
  AO22D0 U103 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), 
        .Z(data_i[5]) );
  AO22D0 U104 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), 
        .Z(data_i[6]) );
  AO22D0 U105 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U106 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U107 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U108 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_15 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AOI221D0 U4 ( .A1(n6), .A2(search_data[31]), .B1(search_data[29]), .B2(n5), 
        .C(n4), .ZN(n19) );
  AOI221D0 U5 ( .A1(n9), .A2(search_data[30]), .B1(search_data[27]), .B2(n8), 
        .C(n7), .ZN(n18) );
  AOI221D0 U6 ( .A1(n12), .A2(search_data[28]), .B1(search_data[24]), .B2(n11), 
        .C(n10), .ZN(n17) );
  AOI221D0 U7 ( .A1(n15), .A2(search_data[26]), .B1(search_data[23]), .B2(n14), 
        .C(n13), .ZN(n16) );
  AOI221D0 U8 ( .A1(n22), .A2(search_data[8]), .B1(search_data[21]), .B2(n21), 
        .C(n20), .ZN(n35) );
  AOI221D0 U9 ( .A1(n25), .A2(search_data[22]), .B1(search_data[19]), .B2(n24), 
        .C(n23), .ZN(n34) );
  AOI221D0 U10 ( .A1(n28), .A2(search_data[20]), .B1(search_data[17]), .B2(n27), .C(n26), .ZN(n33) );
  AOI221D0 U11 ( .A1(n31), .A2(search_data[18]), .B1(search_data[15]), .B2(n30), .C(n29), .ZN(n32) );
  AOI221D0 U12 ( .A1(n38), .A2(search_data[0]), .B1(search_data[13]), .B2(n37), 
        .C(n36), .ZN(n51) );
  AOI221D0 U13 ( .A1(n41), .A2(search_data[14]), .B1(search_data[11]), .B2(n40), .C(n39), .ZN(n50) );
  AOI221D0 U14 ( .A1(n44), .A2(search_data[12]), .B1(search_data[9]), .B2(n43), 
        .C(n42), .ZN(n49) );
  AOI221D0 U15 ( .A1(n47), .A2(search_data[10]), .B1(search_data[25]), .B2(n46), .C(n45), .ZN(n48) );
  AOI221D0 U16 ( .A1(n54), .A2(search_data[7]), .B1(search_data[5]), .B2(n53), 
        .C(n52), .ZN(n65) );
  AOI221D0 U17 ( .A1(n57), .A2(search_data[16]), .B1(search_data[2]), .B2(n56), 
        .C(n55), .ZN(n64) );
  OAI221D0 U18 ( .A1(n60), .A2(search_data[3]), .B1(n59), .B2(search_data[6]), 
        .C(n58), .ZN(n62) );
  CKND0 U19 ( .I(read_value[4]), .ZN(n1) );
  CKND0 U20 ( .I(read_value[1]), .ZN(n2) );
  AOI22D0 U21 ( .A1(search_data[4]), .A2(n1), .B1(search_data[1]), .B2(n2), 
        .ZN(n3) );
  OAI221D0 U22 ( .A1(n1), .A2(search_data[4]), .B1(n2), .B2(search_data[1]), 
        .C(n3), .ZN(n61) );
  AN3D0 U23 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results)
         );
  AO21D0 U24 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U25 ( .A1(reset), .A2(n70), .ZN(n71) );
  CKND2D1 U26 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  AOI21D2 U27 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  CKND0 U28 ( .I(read_value[9]), .ZN(n43) );
  CKND0 U29 ( .I(read_value[10]), .ZN(n47) );
  CKND0 U30 ( .I(read_value[25]), .ZN(n46) );
  CKND0 U31 ( .I(read_value[7]), .ZN(n54) );
  CKND0 U32 ( .I(read_value[12]), .ZN(n44) );
  CKND0 U33 ( .I(read_value[5]), .ZN(n53) );
  CKND0 U34 ( .I(read_value[16]), .ZN(n57) );
  CKND0 U35 ( .I(read_value[2]), .ZN(n56) );
  CKND0 U36 ( .I(read_value[3]), .ZN(n60) );
  CKND0 U37 ( .I(read_value[20]), .ZN(n28) );
  CKND0 U38 ( .I(read_value[17]), .ZN(n27) );
  CKND0 U39 ( .I(read_value[18]), .ZN(n31) );
  CKND0 U40 ( .I(read_value[15]), .ZN(n30) );
  CKND0 U41 ( .I(read_value[0]), .ZN(n38) );
  CKND0 U42 ( .I(read_value[13]), .ZN(n37) );
  CKND0 U43 ( .I(read_value[14]), .ZN(n41) );
  CKND0 U44 ( .I(read_value[11]), .ZN(n40) );
  CKND0 U45 ( .I(read_value[6]), .ZN(n59) );
  CKND0 U46 ( .I(read_value[26]), .ZN(n15) );
  CKND0 U47 ( .I(read_value[24]), .ZN(n11) );
  CKND0 U48 ( .I(read_value[28]), .ZN(n12) );
  CKND0 U49 ( .I(read_value[27]), .ZN(n8) );
  CKND0 U50 ( .I(read_value[23]), .ZN(n14) );
  CKND0 U51 ( .I(read_value[30]), .ZN(n9) );
  CKND0 U52 ( .I(read_value[29]), .ZN(n5) );
  CKND0 U53 ( .I(read_value[31]), .ZN(n6) );
  CKND0 U54 ( .I(read_value[22]), .ZN(n25) );
  CKND0 U55 ( .I(read_value[21]), .ZN(n21) );
  CKND0 U56 ( .I(read_value[8]), .ZN(n22) );
  CKND0 U57 ( .I(read_value[19]), .ZN(n24) );
  AO22D0 U58 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U59 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U60 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U61 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U62 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U63 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U64 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U65 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U66 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U67 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U68 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U69 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U70 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U71 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U72 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U73 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U74 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U75 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U76 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U77 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  ND4D1 U78 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  NR2D1 U79 ( .A1(n62), .A2(n61), .ZN(n63) );
  AOI22D1 U80 ( .A1(search_data[3]), .A2(n60), .B1(search_data[6]), .B2(n59), 
        .ZN(n58) );
  OAI22D1 U81 ( .A1(n57), .A2(search_data[16]), .B1(n56), .B2(search_data[2]), 
        .ZN(n55) );
  OAI22D1 U82 ( .A1(n54), .A2(search_data[7]), .B1(n53), .B2(search_data[5]), 
        .ZN(n52) );
  ND4D1 U83 ( .A1(n51), .A2(n50), .A3(n49), .A4(n48), .ZN(n67) );
  OAI22D1 U84 ( .A1(n47), .A2(search_data[10]), .B1(n46), .B2(search_data[25]), 
        .ZN(n45) );
  OAI22D1 U85 ( .A1(n44), .A2(search_data[12]), .B1(n43), .B2(search_data[9]), 
        .ZN(n42) );
  OAI22D1 U86 ( .A1(n41), .A2(search_data[14]), .B1(n40), .B2(search_data[11]), 
        .ZN(n39) );
  OAI22D1 U87 ( .A1(n38), .A2(search_data[0]), .B1(n37), .B2(search_data[13]), 
        .ZN(n36) );
  ND4D1 U88 ( .A1(n35), .A2(n34), .A3(n33), .A4(n32), .ZN(n68) );
  OAI22D1 U89 ( .A1(n31), .A2(search_data[18]), .B1(n30), .B2(search_data[15]), 
        .ZN(n29) );
  OAI22D1 U90 ( .A1(n28), .A2(search_data[20]), .B1(n27), .B2(search_data[17]), 
        .ZN(n26) );
  OAI22D1 U91 ( .A1(n25), .A2(search_data[22]), .B1(n24), .B2(search_data[19]), 
        .ZN(n23) );
  OAI22D1 U92 ( .A1(n22), .A2(search_data[8]), .B1(n21), .B2(search_data[21]), 
        .ZN(n20) );
  ND4D1 U93 ( .A1(n19), .A2(n18), .A3(n17), .A4(n16), .ZN(n69) );
  OAI22D1 U94 ( .A1(n15), .A2(search_data[26]), .B1(n14), .B2(search_data[23]), 
        .ZN(n13) );
  OAI22D1 U95 ( .A1(n12), .A2(search_data[28]), .B1(n11), .B2(search_data[24]), 
        .ZN(n10) );
  OAI22D1 U96 ( .A1(n9), .A2(search_data[30]), .B1(n8), .B2(search_data[27]), 
        .ZN(n7) );
  OAI22D1 U97 ( .A1(n6), .A2(search_data[31]), .B1(n5), .B2(search_data[29]), 
        .ZN(n4) );
  AO22D0 U98 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U99 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U100 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), 
        .Z(data_i[2]) );
  AO22D0 U101 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), 
        .Z(data_i[3]) );
  AO22D0 U102 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), 
        .Z(data_i[4]) );
  AO22D0 U103 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), 
        .Z(data_i[5]) );
  AO22D0 U104 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), 
        .Z(data_i[6]) );
  AO22D0 U105 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U106 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U107 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U108 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_16 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  OAI22D0 U3 ( .A1(n48), .A2(search_data[19]), .B1(n49), .B2(search_data[22]), 
        .ZN(n1) );
  AOI221D0 U4 ( .A1(n48), .A2(search_data[19]), .B1(search_data[22]), .B2(n49), 
        .C(n1), .ZN(n2) );
  OAI22D0 U5 ( .A1(n46), .A2(search_data[21]), .B1(n47), .B2(search_data[8]), 
        .ZN(n3) );
  AOI221D0 U6 ( .A1(n46), .A2(search_data[21]), .B1(search_data[8]), .B2(n47), 
        .C(n3), .ZN(n4) );
  OAI22D0 U7 ( .A1(n52), .A2(search_data[15]), .B1(n53), .B2(search_data[18]), 
        .ZN(n5) );
  AOI221D0 U8 ( .A1(n52), .A2(search_data[15]), .B1(search_data[18]), .B2(n53), 
        .C(n5), .ZN(n6) );
  OAI22D0 U9 ( .A1(n50), .A2(search_data[17]), .B1(n51), .B2(search_data[20]), 
        .ZN(n7) );
  AOI221D0 U10 ( .A1(n50), .A2(search_data[17]), .B1(search_data[20]), .B2(n51), .C(n7), .ZN(n8) );
  ND4D0 U11 ( .A1(n2), .A2(n4), .A3(n6), .A4(n8), .ZN(n9) );
  OAI22D0 U12 ( .A1(n40), .A2(search_data[27]), .B1(n41), .B2(search_data[30]), 
        .ZN(n10) );
  AOI221D0 U13 ( .A1(n40), .A2(search_data[27]), .B1(search_data[30]), .B2(n41), .C(n10), .ZN(n11) );
  OAI22D0 U14 ( .A1(n38), .A2(search_data[29]), .B1(n39), .B2(search_data[31]), 
        .ZN(n12) );
  AOI221D0 U15 ( .A1(n38), .A2(search_data[29]), .B1(search_data[31]), .B2(n39), .C(n12), .ZN(n13) );
  OAI22D0 U16 ( .A1(n44), .A2(search_data[23]), .B1(n45), .B2(search_data[26]), 
        .ZN(n14) );
  AOI221D0 U17 ( .A1(n44), .A2(search_data[23]), .B1(search_data[26]), .B2(n45), .C(n14), .ZN(n15) );
  OAI22D0 U18 ( .A1(n42), .A2(search_data[24]), .B1(n43), .B2(search_data[28]), 
        .ZN(n16) );
  AOI221D0 U19 ( .A1(n42), .A2(search_data[24]), .B1(search_data[28]), .B2(n43), .C(n16), .ZN(n17) );
  ND4D0 U20 ( .A1(n11), .A2(n13), .A3(n15), .A4(n17), .ZN(n18) );
  AOI22D0 U21 ( .A1(n64), .A2(search_data[7]), .B1(n63), .B2(search_data[5]), 
        .ZN(n19) );
  AO22D0 U22 ( .A1(n67), .A2(search_data[16]), .B1(n66), .B2(search_data[2]), 
        .Z(n20) );
  NR4D0 U23 ( .A1(n65), .A2(n69), .A3(n68), .A4(n20), .ZN(n21) );
  IND4D0 U24 ( .A1(n62), .B1(n19), .B2(search), .B3(n21), .ZN(n22) );
  OAI22D0 U25 ( .A1(n56), .A2(search_data[11]), .B1(n57), .B2(search_data[14]), 
        .ZN(n23) );
  AOI221D0 U26 ( .A1(n56), .A2(search_data[11]), .B1(search_data[14]), .B2(n57), .C(n23), .ZN(n24) );
  OAI22D0 U27 ( .A1(n54), .A2(search_data[13]), .B1(n55), .B2(search_data[0]), 
        .ZN(n25) );
  AOI221D0 U28 ( .A1(n54), .A2(search_data[13]), .B1(search_data[0]), .B2(n55), 
        .C(n25), .ZN(n26) );
  OAI22D0 U29 ( .A1(n60), .A2(search_data[25]), .B1(n61), .B2(search_data[10]), 
        .ZN(n27) );
  AOI221D0 U30 ( .A1(n60), .A2(search_data[25]), .B1(search_data[10]), .B2(n61), .C(n27), .ZN(n28) );
  OAI22D0 U31 ( .A1(n58), .A2(search_data[9]), .B1(n59), .B2(search_data[12]), 
        .ZN(n29) );
  AOI221D0 U32 ( .A1(n58), .A2(search_data[9]), .B1(search_data[12]), .B2(n59), 
        .C(n29), .ZN(n30) );
  ND4D0 U33 ( .A1(n24), .A2(n26), .A3(n28), .A4(n30), .ZN(n31) );
  NR4D0 U34 ( .A1(n9), .A2(n18), .A3(n22), .A4(n31), .ZN(search_results) );
  CKND0 U35 ( .I(read_value[4]), .ZN(n32) );
  CKND0 U36 ( .I(read_value[1]), .ZN(n33) );
  AOI22D0 U37 ( .A1(search_data[4]), .A2(n32), .B1(search_data[1]), .B2(n33), 
        .ZN(n34) );
  OAI221D0 U38 ( .A1(n32), .A2(search_data[4]), .B1(n33), .B2(search_data[1]), 
        .C(n34), .ZN(n68) );
  CKND0 U39 ( .I(read_value[3]), .ZN(n35) );
  CKND0 U40 ( .I(read_value[6]), .ZN(n36) );
  AOI22D0 U41 ( .A1(search_data[6]), .A2(n36), .B1(search_data[3]), .B2(n35), 
        .ZN(n37) );
  OAI221D0 U42 ( .A1(n36), .A2(search_data[6]), .B1(n35), .B2(search_data[3]), 
        .C(n37), .ZN(n69) );
  AN3D0 U43 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results)
         );
  AO21D0 U44 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U45 ( .A1(reset), .A2(n70), .ZN(n71) );
  CKND2D1 U46 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  AOI21D2 U47 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  CKND0 U48 ( .I(read_value[10]), .ZN(n61) );
  CKND0 U49 ( .I(read_value[25]), .ZN(n60) );
  CKND0 U50 ( .I(read_value[18]), .ZN(n53) );
  CKND0 U51 ( .I(read_value[7]), .ZN(n64) );
  CKND0 U52 ( .I(read_value[5]), .ZN(n63) );
  CKND0 U53 ( .I(read_value[0]), .ZN(n55) );
  CKND0 U54 ( .I(read_value[13]), .ZN(n54) );
  CKND0 U55 ( .I(read_value[14]), .ZN(n57) );
  CKND0 U56 ( .I(read_value[11]), .ZN(n56) );
  CKND0 U57 ( .I(read_value[12]), .ZN(n59) );
  CKND0 U58 ( .I(read_value[9]), .ZN(n58) );
  CKND0 U59 ( .I(read_value[15]), .ZN(n52) );
  CKND0 U60 ( .I(read_value[16]), .ZN(n67) );
  CKND0 U61 ( .I(read_value[2]), .ZN(n66) );
  CKND0 U62 ( .I(read_value[23]), .ZN(n44) );
  CKND0 U63 ( .I(read_value[26]), .ZN(n45) );
  CKND0 U64 ( .I(read_value[24]), .ZN(n42) );
  CKND0 U65 ( .I(read_value[28]), .ZN(n43) );
  CKND0 U66 ( .I(read_value[27]), .ZN(n40) );
  CKND0 U67 ( .I(read_value[30]), .ZN(n41) );
  CKND0 U68 ( .I(read_value[31]), .ZN(n39) );
  CKND0 U69 ( .I(read_value[29]), .ZN(n38) );
  CKND0 U70 ( .I(read_value[19]), .ZN(n48) );
  CKND0 U71 ( .I(read_value[22]), .ZN(n49) );
  CKND0 U72 ( .I(read_value[20]), .ZN(n51) );
  CKND0 U73 ( .I(read_value[17]), .ZN(n50) );
  CKND0 U74 ( .I(read_value[8]), .ZN(n47) );
  CKND0 U75 ( .I(read_value[21]), .ZN(n46) );
  AO22D0 U76 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U77 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U78 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), .Z(
        data_i[3]) );
  AO22D0 U79 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U80 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U81 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U82 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), .Z(
        data_i[5]) );
  AO22D0 U83 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U84 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U85 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U86 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U87 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), .Z(
        data_i[2]) );
  AO22D0 U88 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U89 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U90 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U91 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U92 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), .Z(
        data_i[4]) );
  AO22D0 U93 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U94 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), .Z(
        data_i[6]) );
  AO22D0 U95 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  OAI22D1 U96 ( .A1(n67), .A2(search_data[16]), .B1(n66), .B2(search_data[2]), 
        .ZN(n65) );
  OAI22D1 U97 ( .A1(n64), .A2(search_data[7]), .B1(n63), .B2(search_data[5]), 
        .ZN(n62) );
  AO22D0 U98 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U99 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U100 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U101 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U102 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U103 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U104 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U105 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U106 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U107 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U108 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_17 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AOI221D0 U4 ( .A1(n9), .A2(search_data[31]), .B1(search_data[29]), .B2(n8), 
        .C(n7), .ZN(n22) );
  AOI221D0 U5 ( .A1(n12), .A2(search_data[30]), .B1(search_data[27]), .B2(n11), 
        .C(n10), .ZN(n21) );
  AOI221D0 U6 ( .A1(n15), .A2(search_data[28]), .B1(search_data[24]), .B2(n14), 
        .C(n13), .ZN(n20) );
  AOI221D0 U7 ( .A1(n18), .A2(search_data[26]), .B1(search_data[23]), .B2(n17), 
        .C(n16), .ZN(n19) );
  AOI221D0 U8 ( .A1(n25), .A2(search_data[8]), .B1(search_data[21]), .B2(n24), 
        .C(n23), .ZN(n38) );
  AOI221D0 U9 ( .A1(n28), .A2(search_data[22]), .B1(search_data[19]), .B2(n27), 
        .C(n26), .ZN(n37) );
  AOI221D0 U10 ( .A1(n31), .A2(search_data[20]), .B1(search_data[17]), .B2(n30), .C(n29), .ZN(n36) );
  AOI221D0 U11 ( .A1(n34), .A2(search_data[18]), .B1(search_data[15]), .B2(n33), .C(n32), .ZN(n35) );
  AOI221D0 U12 ( .A1(n41), .A2(search_data[0]), .B1(search_data[13]), .B2(n40), 
        .C(n39), .ZN(n54) );
  AOI221D0 U13 ( .A1(n44), .A2(search_data[14]), .B1(search_data[11]), .B2(n43), .C(n42), .ZN(n53) );
  AOI221D0 U14 ( .A1(n47), .A2(search_data[12]), .B1(search_data[9]), .B2(n46), 
        .C(n45), .ZN(n52) );
  AOI221D0 U15 ( .A1(n50), .A2(search_data[10]), .B1(search_data[25]), .B2(n49), .C(n48), .ZN(n51) );
  AOI221D0 U16 ( .A1(n57), .A2(search_data[7]), .B1(search_data[5]), .B2(n56), 
        .C(n55), .ZN(n65) );
  AOI221D0 U17 ( .A1(n60), .A2(search_data[16]), .B1(search_data[2]), .B2(n59), 
        .C(n58), .ZN(n64) );
  CKND0 U18 ( .I(read_value[4]), .ZN(n1) );
  CKND0 U19 ( .I(read_value[1]), .ZN(n2) );
  AOI22D0 U20 ( .A1(search_data[4]), .A2(n1), .B1(search_data[1]), .B2(n2), 
        .ZN(n3) );
  OAI221D0 U21 ( .A1(n1), .A2(search_data[4]), .B1(n2), .B2(search_data[1]), 
        .C(n3), .ZN(n61) );
  CKND0 U22 ( .I(read_value[6]), .ZN(n4) );
  CKND0 U23 ( .I(read_value[3]), .ZN(n5) );
  AOI22D0 U24 ( .A1(search_data[6]), .A2(n4), .B1(search_data[3]), .B2(n5), 
        .ZN(n6) );
  OAI221D0 U25 ( .A1(n4), .A2(search_data[6]), .B1(n5), .B2(search_data[3]), 
        .C(n6), .ZN(n62) );
  AN3D0 U26 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results)
         );
  AO21D0 U27 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U28 ( .A1(reset), .A2(n70), .ZN(n71) );
  CKND2D1 U29 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  AOI21D2 U30 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  OAI22D0 U31 ( .A1(n9), .A2(search_data[31]), .B1(n8), .B2(search_data[29]), 
        .ZN(n7) );
  OAI22D0 U32 ( .A1(n12), .A2(search_data[30]), .B1(n11), .B2(search_data[27]), 
        .ZN(n10) );
  OAI22D0 U33 ( .A1(n34), .A2(search_data[18]), .B1(n33), .B2(search_data[15]), 
        .ZN(n32) );
  OAI22D0 U34 ( .A1(n31), .A2(search_data[20]), .B1(n30), .B2(search_data[17]), 
        .ZN(n29) );
  OAI22D0 U35 ( .A1(n28), .A2(search_data[22]), .B1(n27), .B2(search_data[19]), 
        .ZN(n26) );
  OAI22D0 U36 ( .A1(n41), .A2(search_data[0]), .B1(n40), .B2(search_data[13]), 
        .ZN(n39) );
  OAI22D0 U37 ( .A1(n25), .A2(search_data[8]), .B1(n24), .B2(search_data[21]), 
        .ZN(n23) );
  OAI22D0 U38 ( .A1(n18), .A2(search_data[26]), .B1(n17), .B2(search_data[23]), 
        .ZN(n16) );
  OAI22D0 U39 ( .A1(n15), .A2(search_data[28]), .B1(n14), .B2(search_data[24]), 
        .ZN(n13) );
  OAI22D0 U40 ( .A1(n47), .A2(search_data[12]), .B1(n46), .B2(search_data[9]), 
        .ZN(n45) );
  OAI22D0 U41 ( .A1(n50), .A2(search_data[10]), .B1(n49), .B2(search_data[25]), 
        .ZN(n48) );
  OAI22D0 U42 ( .A1(n60), .A2(search_data[16]), .B1(n59), .B2(search_data[2]), 
        .ZN(n58) );
  OAI22D0 U43 ( .A1(n57), .A2(search_data[7]), .B1(n56), .B2(search_data[5]), 
        .ZN(n55) );
  OAI22D0 U44 ( .A1(n44), .A2(search_data[14]), .B1(n43), .B2(search_data[11]), 
        .ZN(n42) );
  CKND0 U45 ( .I(read_value[16]), .ZN(n60) );
  CKND0 U46 ( .I(read_value[2]), .ZN(n59) );
  CKND0 U47 ( .I(read_value[10]), .ZN(n50) );
  CKND0 U48 ( .I(read_value[25]), .ZN(n49) );
  CKND0 U49 ( .I(read_value[7]), .ZN(n57) );
  CKND0 U50 ( .I(read_value[9]), .ZN(n46) );
  CKND0 U51 ( .I(read_value[5]), .ZN(n56) );
  CKND0 U52 ( .I(read_value[12]), .ZN(n47) );
  CKND0 U53 ( .I(read_value[8]), .ZN(n25) );
  CKND0 U54 ( .I(read_value[18]), .ZN(n34) );
  CKND0 U55 ( .I(read_value[31]), .ZN(n9) );
  CKND0 U56 ( .I(read_value[29]), .ZN(n8) );
  CKND0 U57 ( .I(read_value[17]), .ZN(n30) );
  CKND0 U58 ( .I(read_value[30]), .ZN(n12) );
  CKND0 U59 ( .I(read_value[27]), .ZN(n11) );
  CKND0 U60 ( .I(read_value[20]), .ZN(n31) );
  CKND0 U61 ( .I(read_value[28]), .ZN(n15) );
  CKND0 U62 ( .I(read_value[24]), .ZN(n14) );
  CKND0 U63 ( .I(read_value[19]), .ZN(n27) );
  CKND0 U64 ( .I(read_value[26]), .ZN(n18) );
  CKND0 U65 ( .I(read_value[23]), .ZN(n17) );
  CKND0 U66 ( .I(read_value[21]), .ZN(n24) );
  CKND0 U67 ( .I(read_value[13]), .ZN(n40) );
  CKND0 U68 ( .I(read_value[0]), .ZN(n41) );
  CKND0 U69 ( .I(read_value[14]), .ZN(n44) );
  CKND0 U70 ( .I(read_value[15]), .ZN(n33) );
  CKND0 U71 ( .I(read_value[22]), .ZN(n28) );
  CKND0 U72 ( .I(read_value[11]), .ZN(n43) );
  AO22D0 U73 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U74 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U75 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U76 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U77 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), .Z(
        data_i[6]) );
  AO22D0 U78 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U79 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), .Z(
        data_i[5]) );
  AO22D0 U80 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U81 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), .Z(
        data_i[4]) );
  AO22D0 U82 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), .Z(
        data_i[3]) );
  AO22D0 U83 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), .Z(
        data_i[2]) );
  AO22D0 U84 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U85 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U86 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U87 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U88 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U89 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U90 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U91 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U92 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  ND4D1 U93 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  NR2D1 U94 ( .A1(n62), .A2(n61), .ZN(n63) );
  ND4D1 U95 ( .A1(n54), .A2(n53), .A3(n52), .A4(n51), .ZN(n67) );
  ND4D1 U96 ( .A1(n38), .A2(n37), .A3(n36), .A4(n35), .ZN(n68) );
  ND4D1 U97 ( .A1(n22), .A2(n21), .A3(n20), .A4(n19), .ZN(n69) );
  AO22D0 U98 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U99 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U100 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U101 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U102 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U103 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U104 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U105 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U106 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U107 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U108 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_18 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  CKND0 U3 ( .I(read_value[4]), .ZN(n1) );
  CKND0 U4 ( .I(read_value[1]), .ZN(n2) );
  AOI22D0 U5 ( .A1(search_data[4]), .A2(n1), .B1(search_data[1]), .B2(n2), 
        .ZN(n3) );
  OAI221D0 U6 ( .A1(n1), .A2(search_data[4]), .B1(n2), .B2(search_data[1]), 
        .C(n3), .ZN(n68) );
  OAI22D0 U7 ( .A1(n46), .A2(search_data[19]), .B1(n47), .B2(search_data[22]), 
        .ZN(n4) );
  AOI221D0 U8 ( .A1(n46), .A2(search_data[19]), .B1(search_data[22]), .B2(n47), 
        .C(n4), .ZN(n5) );
  OAI22D0 U9 ( .A1(n44), .A2(search_data[21]), .B1(n45), .B2(search_data[8]), 
        .ZN(n6) );
  AOI221D0 U10 ( .A1(n44), .A2(search_data[21]), .B1(search_data[8]), .B2(n45), 
        .C(n6), .ZN(n7) );
  OAI22D0 U11 ( .A1(n50), .A2(search_data[15]), .B1(n51), .B2(search_data[18]), 
        .ZN(n8) );
  AOI221D0 U12 ( .A1(n50), .A2(search_data[15]), .B1(search_data[18]), .B2(n51), .C(n8), .ZN(n9) );
  OAI22D0 U13 ( .A1(n48), .A2(search_data[17]), .B1(n49), .B2(search_data[20]), 
        .ZN(n10) );
  AOI221D0 U14 ( .A1(n48), .A2(search_data[17]), .B1(search_data[20]), .B2(n49), .C(n10), .ZN(n11) );
  ND4D0 U15 ( .A1(n5), .A2(n7), .A3(n9), .A4(n11), .ZN(n12) );
  OAI22D0 U16 ( .A1(n38), .A2(search_data[27]), .B1(n39), .B2(search_data[30]), 
        .ZN(n13) );
  AOI221D0 U17 ( .A1(n38), .A2(search_data[27]), .B1(search_data[30]), .B2(n39), .C(n13), .ZN(n14) );
  OAI22D0 U18 ( .A1(n36), .A2(search_data[29]), .B1(n37), .B2(search_data[31]), 
        .ZN(n15) );
  AOI221D0 U19 ( .A1(n36), .A2(search_data[29]), .B1(search_data[31]), .B2(n37), .C(n15), .ZN(n16) );
  OAI22D0 U20 ( .A1(n42), .A2(search_data[23]), .B1(n43), .B2(search_data[26]), 
        .ZN(n17) );
  AOI221D0 U21 ( .A1(n42), .A2(search_data[23]), .B1(search_data[26]), .B2(n43), .C(n17), .ZN(n18) );
  OAI22D0 U22 ( .A1(n40), .A2(search_data[24]), .B1(n41), .B2(search_data[28]), 
        .ZN(n19) );
  AOI221D0 U23 ( .A1(n40), .A2(search_data[24]), .B1(search_data[28]), .B2(n41), .C(n19), .ZN(n20) );
  ND4D0 U24 ( .A1(n14), .A2(n16), .A3(n18), .A4(n20), .ZN(n21) );
  OAI22D0 U25 ( .A1(n60), .A2(search_data[5]), .B1(n61), .B2(search_data[7]), 
        .ZN(n22) );
  AOI221D0 U26 ( .A1(n60), .A2(search_data[5]), .B1(search_data[7]), .B2(n61), 
        .C(n22), .ZN(n23) );
  AO22D0 U27 ( .A1(n64), .A2(search_data[16]), .B1(n63), .B2(search_data[2]), 
        .Z(n24) );
  NR4D0 U28 ( .A1(n62), .A2(n69), .A3(n68), .A4(n24), .ZN(n25) );
  AOI22D0 U29 ( .A1(n55), .A2(search_data[14]), .B1(n54), .B2(search_data[11]), 
        .ZN(n26) );
  OAI221D0 U30 ( .A1(n55), .A2(search_data[14]), .B1(n54), .B2(search_data[11]), .C(n26), .ZN(n27) );
  AOI22D0 U31 ( .A1(n53), .A2(search_data[0]), .B1(n52), .B2(search_data[13]), 
        .ZN(n28) );
  OAI221D0 U32 ( .A1(n53), .A2(search_data[0]), .B1(n52), .B2(search_data[13]), 
        .C(n28), .ZN(n29) );
  AOI22D0 U33 ( .A1(n59), .A2(search_data[10]), .B1(n58), .B2(search_data[25]), 
        .ZN(n30) );
  OAI221D0 U34 ( .A1(n59), .A2(search_data[10]), .B1(n58), .B2(search_data[25]), .C(n30), .ZN(n31) );
  AOI22D0 U35 ( .A1(n57), .A2(search_data[12]), .B1(n56), .B2(search_data[9]), 
        .ZN(n32) );
  OAI221D0 U36 ( .A1(n57), .A2(search_data[12]), .B1(n56), .B2(search_data[9]), 
        .C(n32), .ZN(n33) );
  NR4D0 U37 ( .A1(n27), .A2(n29), .A3(n31), .A4(n33), .ZN(n34) );
  ND4D0 U38 ( .A1(n23), .A2(search), .A3(n25), .A4(n34), .ZN(n35) );
  NR3D0 U39 ( .A1(n12), .A2(n21), .A3(n35), .ZN(search_results) );
  AN3D0 U40 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results)
         );
  AO21D0 U41 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U42 ( .A1(reset), .A2(n70), .ZN(n71) );
  CKND2D1 U43 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  AOI21D2 U44 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  OAI22D0 U45 ( .A1(n64), .A2(search_data[16]), .B1(n63), .B2(search_data[2]), 
        .ZN(n62) );
  AOI22D0 U46 ( .A1(search_data[3]), .A2(n67), .B1(search_data[6]), .B2(n66), 
        .ZN(n65) );
  CKND0 U47 ( .I(read_value[10]), .ZN(n59) );
  CKND0 U48 ( .I(read_value[13]), .ZN(n52) );
  CKND0 U49 ( .I(read_value[12]), .ZN(n57) );
  CKND0 U50 ( .I(read_value[0]), .ZN(n53) );
  CKND0 U51 ( .I(read_value[25]), .ZN(n58) );
  CKND0 U52 ( .I(read_value[9]), .ZN(n56) );
  CKND0 U53 ( .I(read_value[11]), .ZN(n54) );
  CKND0 U54 ( .I(read_value[14]), .ZN(n55) );
  CKND0 U55 ( .I(read_value[27]), .ZN(n38) );
  CKND0 U56 ( .I(read_value[20]), .ZN(n49) );
  CKND0 U57 ( .I(read_value[28]), .ZN(n41) );
  CKND0 U58 ( .I(read_value[24]), .ZN(n40) );
  CKND0 U59 ( .I(read_value[19]), .ZN(n46) );
  CKND0 U60 ( .I(read_value[16]), .ZN(n64) );
  CKND0 U61 ( .I(read_value[26]), .ZN(n43) );
  CKND0 U62 ( .I(read_value[6]), .ZN(n66) );
  CKND0 U63 ( .I(read_value[23]), .ZN(n42) );
  CKND0 U64 ( .I(read_value[3]), .ZN(n67) );
  CKND0 U65 ( .I(read_value[22]), .ZN(n47) );
  CKND0 U66 ( .I(read_value[2]), .ZN(n63) );
  CKND0 U67 ( .I(read_value[8]), .ZN(n45) );
  CKND0 U68 ( .I(read_value[21]), .ZN(n44) );
  CKND0 U69 ( .I(read_value[15]), .ZN(n50) );
  CKND0 U70 ( .I(read_value[18]), .ZN(n51) );
  CKND0 U71 ( .I(read_value[7]), .ZN(n61) );
  CKND0 U72 ( .I(read_value[31]), .ZN(n37) );
  CKND0 U73 ( .I(read_value[29]), .ZN(n36) );
  CKND0 U74 ( .I(read_value[17]), .ZN(n48) );
  CKND0 U75 ( .I(read_value[5]), .ZN(n60) );
  CKND0 U76 ( .I(read_value[30]), .ZN(n39) );
  AO22D0 U77 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U78 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U79 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), .Z(
        data_i[3]) );
  AO22D0 U80 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), .Z(
        data_i[4]) );
  AO22D0 U81 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), .Z(
        data_i[5]) );
  AO22D0 U82 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), .Z(
        data_i[6]) );
  AO22D0 U83 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U84 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U85 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), .Z(
        data_i[2]) );
  AO22D0 U86 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U87 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U88 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U89 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U90 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U91 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U92 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U93 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U94 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U95 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U96 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  OAI221D0 U97 ( .A1(n67), .A2(search_data[3]), .B1(n66), .B2(search_data[6]), 
        .C(n65), .ZN(n69) );
  AO22D0 U98 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U99 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U100 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U101 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U102 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U103 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U104 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U105 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U106 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U107 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U108 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_19 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AN3D0 U4 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results) );
  AO21D0 U5 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U6 ( .A1(reset), .A2(n70), .ZN(n71) );
  CKND2D1 U7 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  AOI21D2 U8 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  OAI22D0 U9 ( .A1(n44), .A2(search_data[10]), .B1(n43), .B2(search_data[25]), 
        .ZN(n42) );
  OAI22D0 U10 ( .A1(n19), .A2(search_data[8]), .B1(n18), .B2(search_data[21]), 
        .ZN(n17) );
  OAI22D0 U11 ( .A1(n51), .A2(search_data[7]), .B1(n50), .B2(search_data[5]), 
        .ZN(n49) );
  OAI22D0 U12 ( .A1(n12), .A2(search_data[26]), .B1(n11), .B2(search_data[23]), 
        .ZN(n10) );
  OAI22D0 U13 ( .A1(n54), .A2(search_data[16]), .B1(n53), .B2(search_data[2]), 
        .ZN(n52) );
  OAI22D0 U14 ( .A1(n9), .A2(search_data[28]), .B1(n8), .B2(search_data[24]), 
        .ZN(n7) );
  AOI22D0 U15 ( .A1(search_data[3]), .A2(n57), .B1(search_data[6]), .B2(n56), 
        .ZN(n55) );
  OAI22D0 U16 ( .A1(n6), .A2(search_data[30]), .B1(n5), .B2(search_data[27]), 
        .ZN(n4) );
  AOI22D0 U17 ( .A1(search_data[1]), .A2(n60), .B1(search_data[4]), .B2(n59), 
        .ZN(n58) );
  OAI22D0 U18 ( .A1(n3), .A2(search_data[31]), .B1(n2), .B2(search_data[29]), 
        .ZN(n1) );
  OAI22D0 U19 ( .A1(n28), .A2(search_data[18]), .B1(n27), .B2(search_data[15]), 
        .ZN(n26) );
  OAI22D0 U20 ( .A1(n35), .A2(search_data[0]), .B1(n34), .B2(search_data[13]), 
        .ZN(n33) );
  OAI22D0 U21 ( .A1(n25), .A2(search_data[20]), .B1(n24), .B2(search_data[17]), 
        .ZN(n23) );
  OAI22D0 U22 ( .A1(n38), .A2(search_data[14]), .B1(n37), .B2(search_data[11]), 
        .ZN(n36) );
  OAI22D0 U23 ( .A1(n22), .A2(search_data[22]), .B1(n21), .B2(search_data[19]), 
        .ZN(n20) );
  OAI22D0 U24 ( .A1(n41), .A2(search_data[12]), .B1(n40), .B2(search_data[9]), 
        .ZN(n39) );
  CKND0 U25 ( .I(read_value[13]), .ZN(n34) );
  CKND0 U26 ( .I(read_value[22]), .ZN(n22) );
  CKND0 U27 ( .I(read_value[14]), .ZN(n38) );
  CKND0 U28 ( .I(read_value[11]), .ZN(n37) );
  CKND0 U29 ( .I(read_value[24]), .ZN(n8) );
  CKND0 U30 ( .I(read_value[21]), .ZN(n18) );
  CKND0 U31 ( .I(read_value[12]), .ZN(n41) );
  CKND0 U32 ( .I(read_value[20]), .ZN(n25) );
  CKND0 U33 ( .I(read_value[17]), .ZN(n24) );
  CKND0 U34 ( .I(read_value[8]), .ZN(n19) );
  CKND0 U35 ( .I(read_value[18]), .ZN(n28) );
  CKND0 U36 ( .I(read_value[19]), .ZN(n21) );
  CKND0 U37 ( .I(read_value[23]), .ZN(n11) );
  CKND0 U38 ( .I(read_value[15]), .ZN(n27) );
  CKND0 U39 ( .I(read_value[0]), .ZN(n35) );
  CKND0 U40 ( .I(read_value[26]), .ZN(n12) );
  CKND0 U41 ( .I(read_value[3]), .ZN(n57) );
  CKND0 U42 ( .I(read_value[6]), .ZN(n56) );
  CKND0 U43 ( .I(read_value[1]), .ZN(n60) );
  CKND0 U44 ( .I(read_value[4]), .ZN(n59) );
  CKND0 U45 ( .I(read_value[9]), .ZN(n40) );
  CKND0 U46 ( .I(read_value[28]), .ZN(n9) );
  CKND0 U47 ( .I(read_value[27]), .ZN(n5) );
  CKND0 U48 ( .I(read_value[10]), .ZN(n44) );
  CKND0 U49 ( .I(read_value[25]), .ZN(n43) );
  CKND0 U50 ( .I(read_value[30]), .ZN(n6) );
  CKND0 U51 ( .I(read_value[7]), .ZN(n51) );
  CKND0 U52 ( .I(read_value[5]), .ZN(n50) );
  CKND0 U53 ( .I(read_value[29]), .ZN(n2) );
  CKND0 U54 ( .I(read_value[16]), .ZN(n54) );
  CKND0 U55 ( .I(read_value[31]), .ZN(n3) );
  CKND0 U56 ( .I(read_value[2]), .ZN(n53) );
  AO22D0 U57 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U58 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U59 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U60 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), .Z(
        data_i[2]) );
  AO22D0 U61 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), .Z(
        data_i[3]) );
  AO22D0 U62 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), .Z(
        data_i[4]) );
  AO22D0 U63 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), .Z(
        data_i[5]) );
  AO22D0 U64 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), .Z(
        data_i[6]) );
  AO22D0 U65 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U66 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U67 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U68 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U69 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U70 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U71 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U72 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U73 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U74 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U75 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U76 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  ND4D1 U77 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  NR2D1 U78 ( .A1(n62), .A2(n61), .ZN(n63) );
  ND4D1 U79 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .ZN(n67) );
  ND4D1 U80 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .ZN(n68) );
  ND4D1 U81 ( .A1(n16), .A2(n15), .A3(n14), .A4(n13), .ZN(n69) );
  AOI221D0 U82 ( .A1(n3), .A2(search_data[31]), .B1(search_data[29]), .B2(n2), 
        .C(n1), .ZN(n16) );
  AOI221D0 U83 ( .A1(n6), .A2(search_data[30]), .B1(search_data[27]), .B2(n5), 
        .C(n4), .ZN(n15) );
  AOI221D0 U84 ( .A1(n9), .A2(search_data[28]), .B1(search_data[24]), .B2(n8), 
        .C(n7), .ZN(n14) );
  AOI221D0 U85 ( .A1(n12), .A2(search_data[26]), .B1(search_data[23]), .B2(n11), .C(n10), .ZN(n13) );
  AOI221D0 U86 ( .A1(n19), .A2(search_data[8]), .B1(search_data[21]), .B2(n18), 
        .C(n17), .ZN(n32) );
  AOI221D0 U87 ( .A1(n22), .A2(search_data[22]), .B1(search_data[19]), .B2(n21), .C(n20), .ZN(n31) );
  AOI221D0 U88 ( .A1(n25), .A2(search_data[20]), .B1(search_data[17]), .B2(n24), .C(n23), .ZN(n30) );
  AOI221D0 U89 ( .A1(n28), .A2(search_data[18]), .B1(search_data[15]), .B2(n27), .C(n26), .ZN(n29) );
  AOI221D0 U90 ( .A1(n35), .A2(search_data[0]), .B1(search_data[13]), .B2(n34), 
        .C(n33), .ZN(n48) );
  AOI221D0 U91 ( .A1(n38), .A2(search_data[14]), .B1(search_data[11]), .B2(n37), .C(n36), .ZN(n47) );
  AOI221D0 U92 ( .A1(n41), .A2(search_data[12]), .B1(search_data[9]), .B2(n40), 
        .C(n39), .ZN(n46) );
  AOI221D0 U93 ( .A1(n44), .A2(search_data[10]), .B1(search_data[25]), .B2(n43), .C(n42), .ZN(n45) );
  AOI221D0 U94 ( .A1(n51), .A2(search_data[7]), .B1(search_data[5]), .B2(n50), 
        .C(n49), .ZN(n65) );
  AOI221D0 U95 ( .A1(n54), .A2(search_data[16]), .B1(search_data[2]), .B2(n53), 
        .C(n52), .ZN(n64) );
  OAI221D0 U96 ( .A1(n57), .A2(search_data[3]), .B1(n56), .B2(search_data[6]), 
        .C(n55), .ZN(n62) );
  OAI221D0 U97 ( .A1(n60), .A2(search_data[1]), .B1(n59), .B2(search_data[4]), 
        .C(n58), .ZN(n61) );
  AO22D0 U98 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U99 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U100 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U101 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U102 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U103 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U104 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U105 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U106 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U107 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U108 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_20 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AN3D0 U4 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results) );
  ND4D0 U5 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  AO21D0 U6 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U7 ( .A1(reset), .A2(n70), .ZN(n71) );
  CKND2D1 U8 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  AOI21D2 U9 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  AOI22D0 U10 ( .A1(search_data[1]), .A2(n60), .B1(search_data[4]), .B2(n59), 
        .ZN(n58) );
  OAI22D0 U11 ( .A1(n38), .A2(search_data[14]), .B1(n37), .B2(search_data[11]), 
        .ZN(n36) );
  OAI22D0 U12 ( .A1(n35), .A2(search_data[0]), .B1(n34), .B2(search_data[13]), 
        .ZN(n33) );
  OAI22D0 U13 ( .A1(n28), .A2(search_data[18]), .B1(n27), .B2(search_data[15]), 
        .ZN(n26) );
  OAI22D0 U14 ( .A1(n25), .A2(search_data[20]), .B1(n24), .B2(search_data[17]), 
        .ZN(n23) );
  OAI22D0 U15 ( .A1(n22), .A2(search_data[22]), .B1(n21), .B2(search_data[19]), 
        .ZN(n20) );
  OAI22D0 U16 ( .A1(n19), .A2(search_data[8]), .B1(n18), .B2(search_data[21]), 
        .ZN(n17) );
  OAI22D0 U17 ( .A1(n12), .A2(search_data[26]), .B1(n11), .B2(search_data[23]), 
        .ZN(n10) );
  OAI22D0 U18 ( .A1(n9), .A2(search_data[28]), .B1(n8), .B2(search_data[24]), 
        .ZN(n7) );
  OAI22D0 U19 ( .A1(n6), .A2(search_data[30]), .B1(n5), .B2(search_data[27]), 
        .ZN(n4) );
  AOI22D0 U20 ( .A1(search_data[3]), .A2(n57), .B1(search_data[6]), .B2(n56), 
        .ZN(n55) );
  OAI22D0 U21 ( .A1(n54), .A2(search_data[16]), .B1(n53), .B2(search_data[2]), 
        .ZN(n52) );
  OAI22D0 U22 ( .A1(n51), .A2(search_data[7]), .B1(n50), .B2(search_data[5]), 
        .ZN(n49) );
  OAI22D0 U23 ( .A1(n44), .A2(search_data[10]), .B1(n43), .B2(search_data[25]), 
        .ZN(n42) );
  OAI22D0 U24 ( .A1(n3), .A2(search_data[31]), .B1(n2), .B2(search_data[29]), 
        .ZN(n1) );
  OAI22D0 U25 ( .A1(n41), .A2(search_data[12]), .B1(n40), .B2(search_data[9]), 
        .ZN(n39) );
  CKND0 U26 ( .I(read_value[13]), .ZN(n34) );
  CKND0 U27 ( .I(read_value[15]), .ZN(n27) );
  CKND0 U28 ( .I(read_value[10]), .ZN(n44) );
  CKND0 U29 ( .I(read_value[0]), .ZN(n35) );
  CKND0 U30 ( .I(read_value[25]), .ZN(n43) );
  CKND0 U31 ( .I(read_value[19]), .ZN(n21) );
  CKND0 U32 ( .I(read_value[22]), .ZN(n22) );
  CKND0 U33 ( .I(read_value[18]), .ZN(n28) );
  CKND0 U34 ( .I(read_value[14]), .ZN(n38) );
  CKND0 U35 ( .I(read_value[11]), .ZN(n37) );
  CKND0 U36 ( .I(read_value[12]), .ZN(n41) );
  CKND0 U37 ( .I(read_value[17]), .ZN(n24) );
  CKND0 U38 ( .I(read_value[9]), .ZN(n40) );
  CKND0 U39 ( .I(read_value[20]), .ZN(n25) );
  CKND0 U40 ( .I(read_value[26]), .ZN(n12) );
  CKND0 U41 ( .I(read_value[1]), .ZN(n60) );
  CKND0 U42 ( .I(read_value[4]), .ZN(n59) );
  CKND0 U43 ( .I(read_value[24]), .ZN(n8) );
  CKND0 U44 ( .I(read_value[31]), .ZN(n3) );
  CKND0 U45 ( .I(read_value[29]), .ZN(n2) );
  CKND0 U46 ( .I(read_value[28]), .ZN(n9) );
  CKND0 U47 ( .I(read_value[30]), .ZN(n6) );
  CKND0 U48 ( .I(read_value[27]), .ZN(n5) );
  CKND0 U49 ( .I(read_value[7]), .ZN(n51) );
  CKND0 U50 ( .I(read_value[5]), .ZN(n50) );
  CKND0 U51 ( .I(read_value[16]), .ZN(n54) );
  CKND0 U52 ( .I(read_value[21]), .ZN(n18) );
  CKND0 U53 ( .I(read_value[2]), .ZN(n53) );
  CKND0 U54 ( .I(read_value[8]), .ZN(n19) );
  CKND0 U55 ( .I(read_value[3]), .ZN(n57) );
  CKND0 U56 ( .I(read_value[6]), .ZN(n56) );
  CKND0 U57 ( .I(read_value[23]), .ZN(n11) );
  AO22D0 U58 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U59 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), .Z(
        data_i[3]) );
  AO22D0 U60 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), .Z(
        data_i[4]) );
  AO22D0 U61 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U62 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U63 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), .Z(
        data_i[6]) );
  AO22D0 U64 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), .Z(
        data_i[2]) );
  AO22D0 U65 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U66 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U67 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U68 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U69 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U70 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U71 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), .Z(
        data_i[5]) );
  AO22D0 U72 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U73 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U74 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U75 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U76 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U77 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  NR2D1 U78 ( .A1(n62), .A2(n61), .ZN(n63) );
  ND4D1 U79 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .ZN(n67) );
  ND4D1 U80 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .ZN(n68) );
  ND4D1 U81 ( .A1(n16), .A2(n15), .A3(n14), .A4(n13), .ZN(n69) );
  AOI221D0 U82 ( .A1(n3), .A2(search_data[31]), .B1(search_data[29]), .B2(n2), 
        .C(n1), .ZN(n16) );
  AOI221D0 U83 ( .A1(n6), .A2(search_data[30]), .B1(search_data[27]), .B2(n5), 
        .C(n4), .ZN(n15) );
  AOI221D0 U84 ( .A1(n9), .A2(search_data[28]), .B1(search_data[24]), .B2(n8), 
        .C(n7), .ZN(n14) );
  AOI221D0 U85 ( .A1(n12), .A2(search_data[26]), .B1(search_data[23]), .B2(n11), .C(n10), .ZN(n13) );
  AOI221D0 U86 ( .A1(n19), .A2(search_data[8]), .B1(search_data[21]), .B2(n18), 
        .C(n17), .ZN(n32) );
  AOI221D0 U87 ( .A1(n22), .A2(search_data[22]), .B1(search_data[19]), .B2(n21), .C(n20), .ZN(n31) );
  AOI221D0 U88 ( .A1(n25), .A2(search_data[20]), .B1(search_data[17]), .B2(n24), .C(n23), .ZN(n30) );
  AOI221D0 U89 ( .A1(n28), .A2(search_data[18]), .B1(search_data[15]), .B2(n27), .C(n26), .ZN(n29) );
  AOI221D0 U90 ( .A1(n35), .A2(search_data[0]), .B1(search_data[13]), .B2(n34), 
        .C(n33), .ZN(n48) );
  AOI221D0 U91 ( .A1(n38), .A2(search_data[14]), .B1(search_data[11]), .B2(n37), .C(n36), .ZN(n47) );
  AOI221D0 U92 ( .A1(n41), .A2(search_data[12]), .B1(search_data[9]), .B2(n40), 
        .C(n39), .ZN(n46) );
  AOI221D0 U93 ( .A1(n44), .A2(search_data[10]), .B1(search_data[25]), .B2(n43), .C(n42), .ZN(n45) );
  AOI221D0 U94 ( .A1(n51), .A2(search_data[7]), .B1(search_data[5]), .B2(n50), 
        .C(n49), .ZN(n65) );
  AOI221D0 U95 ( .A1(n54), .A2(search_data[16]), .B1(search_data[2]), .B2(n53), 
        .C(n52), .ZN(n64) );
  OAI221D0 U96 ( .A1(n57), .A2(search_data[3]), .B1(n56), .B2(search_data[6]), 
        .C(n55), .ZN(n62) );
  OAI221D0 U97 ( .A1(n60), .A2(search_data[1]), .B1(n59), .B2(search_data[4]), 
        .C(n58), .ZN(n61) );
  AO22D0 U98 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U99 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U100 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U101 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U102 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U103 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U104 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U105 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U106 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U107 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U108 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_21 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AN3D0 U4 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results) );
  ND4D0 U5 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  AO21D0 U6 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U7 ( .A1(reset), .A2(n70), .ZN(n71) );
  CKND2D1 U8 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  AOI21D2 U9 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  OAI22D0 U10 ( .A1(n3), .A2(search_data[31]), .B1(n2), .B2(search_data[29]), 
        .ZN(n1) );
  OAI22D0 U11 ( .A1(n6), .A2(search_data[30]), .B1(n5), .B2(search_data[27]), 
        .ZN(n4) );
  OAI22D0 U12 ( .A1(n9), .A2(search_data[28]), .B1(n8), .B2(search_data[24]), 
        .ZN(n7) );
  OAI22D0 U13 ( .A1(n12), .A2(search_data[26]), .B1(n11), .B2(search_data[23]), 
        .ZN(n10) );
  OAI22D0 U14 ( .A1(n19), .A2(search_data[8]), .B1(n18), .B2(search_data[21]), 
        .ZN(n17) );
  OAI22D0 U15 ( .A1(n22), .A2(search_data[22]), .B1(n21), .B2(search_data[19]), 
        .ZN(n20) );
  OAI22D0 U16 ( .A1(n25), .A2(search_data[20]), .B1(n24), .B2(search_data[17]), 
        .ZN(n23) );
  OAI22D0 U17 ( .A1(n28), .A2(search_data[18]), .B1(n27), .B2(search_data[15]), 
        .ZN(n26) );
  OAI22D0 U18 ( .A1(n35), .A2(search_data[0]), .B1(n34), .B2(search_data[13]), 
        .ZN(n33) );
  OAI22D0 U19 ( .A1(n38), .A2(search_data[14]), .B1(n37), .B2(search_data[11]), 
        .ZN(n36) );
  OAI22D0 U20 ( .A1(n41), .A2(search_data[12]), .B1(n40), .B2(search_data[9]), 
        .ZN(n39) );
  OAI22D0 U21 ( .A1(n44), .A2(search_data[10]), .B1(n43), .B2(search_data[25]), 
        .ZN(n42) );
  OAI22D0 U22 ( .A1(n51), .A2(search_data[7]), .B1(n50), .B2(search_data[5]), 
        .ZN(n49) );
  OAI22D0 U23 ( .A1(n54), .A2(search_data[16]), .B1(n53), .B2(search_data[2]), 
        .ZN(n52) );
  AOI22D0 U24 ( .A1(search_data[3]), .A2(n57), .B1(search_data[6]), .B2(n56), 
        .ZN(n55) );
  AOI22D0 U25 ( .A1(search_data[1]), .A2(n60), .B1(search_data[4]), .B2(n59), 
        .ZN(n58) );
  CKND0 U26 ( .I(read_value[1]), .ZN(n60) );
  CKND0 U27 ( .I(read_value[4]), .ZN(n59) );
  CKND0 U28 ( .I(read_value[6]), .ZN(n56) );
  CKND0 U29 ( .I(read_value[3]), .ZN(n57) );
  CKND0 U30 ( .I(read_value[2]), .ZN(n53) );
  CKND0 U31 ( .I(read_value[16]), .ZN(n54) );
  CKND0 U32 ( .I(read_value[18]), .ZN(n28) );
  CKND0 U33 ( .I(read_value[17]), .ZN(n24) );
  CKND0 U34 ( .I(read_value[20]), .ZN(n25) );
  CKND0 U35 ( .I(read_value[19]), .ZN(n21) );
  CKND0 U36 ( .I(read_value[22]), .ZN(n22) );
  CKND0 U37 ( .I(read_value[21]), .ZN(n18) );
  CKND0 U38 ( .I(read_value[8]), .ZN(n19) );
  CKND0 U39 ( .I(read_value[31]), .ZN(n3) );
  CKND0 U40 ( .I(read_value[23]), .ZN(n11) );
  CKND0 U41 ( .I(read_value[26]), .ZN(n12) );
  CKND0 U42 ( .I(read_value[29]), .ZN(n2) );
  CKND0 U43 ( .I(read_value[24]), .ZN(n8) );
  CKND0 U44 ( .I(read_value[28]), .ZN(n9) );
  CKND0 U45 ( .I(read_value[27]), .ZN(n5) );
  CKND0 U46 ( .I(read_value[15]), .ZN(n27) );
  CKND0 U47 ( .I(read_value[5]), .ZN(n50) );
  CKND0 U48 ( .I(read_value[7]), .ZN(n51) );
  CKND0 U49 ( .I(read_value[25]), .ZN(n43) );
  CKND0 U50 ( .I(read_value[10]), .ZN(n44) );
  CKND0 U51 ( .I(read_value[9]), .ZN(n40) );
  CKND0 U52 ( .I(read_value[12]), .ZN(n41) );
  CKND0 U53 ( .I(read_value[11]), .ZN(n37) );
  CKND0 U54 ( .I(read_value[14]), .ZN(n38) );
  CKND0 U55 ( .I(read_value[13]), .ZN(n34) );
  CKND0 U56 ( .I(read_value[0]), .ZN(n35) );
  CKND0 U57 ( .I(read_value[30]), .ZN(n6) );
  AO22D0 U58 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U59 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U60 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), .Z(
        data_i[2]) );
  AO22D0 U61 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), .Z(
        data_i[3]) );
  AO22D0 U62 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), .Z(
        data_i[4]) );
  AO22D0 U63 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), .Z(
        data_i[5]) );
  AO22D0 U64 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), .Z(
        data_i[6]) );
  AO22D0 U65 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U66 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U67 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U68 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U69 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U70 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U71 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U72 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U73 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U74 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U75 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U76 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U77 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  NR2D1 U78 ( .A1(n62), .A2(n61), .ZN(n63) );
  ND4D1 U79 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .ZN(n67) );
  ND4D1 U80 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .ZN(n68) );
  ND4D1 U81 ( .A1(n16), .A2(n15), .A3(n14), .A4(n13), .ZN(n69) );
  AOI221D0 U82 ( .A1(n3), .A2(search_data[31]), .B1(search_data[29]), .B2(n2), 
        .C(n1), .ZN(n16) );
  AOI221D0 U83 ( .A1(n6), .A2(search_data[30]), .B1(search_data[27]), .B2(n5), 
        .C(n4), .ZN(n15) );
  AOI221D0 U84 ( .A1(n9), .A2(search_data[28]), .B1(search_data[24]), .B2(n8), 
        .C(n7), .ZN(n14) );
  AOI221D0 U85 ( .A1(n12), .A2(search_data[26]), .B1(search_data[23]), .B2(n11), .C(n10), .ZN(n13) );
  AOI221D0 U86 ( .A1(n19), .A2(search_data[8]), .B1(search_data[21]), .B2(n18), 
        .C(n17), .ZN(n32) );
  AOI221D0 U87 ( .A1(n22), .A2(search_data[22]), .B1(search_data[19]), .B2(n21), .C(n20), .ZN(n31) );
  AOI221D0 U88 ( .A1(n25), .A2(search_data[20]), .B1(search_data[17]), .B2(n24), .C(n23), .ZN(n30) );
  AOI221D0 U89 ( .A1(n28), .A2(search_data[18]), .B1(search_data[15]), .B2(n27), .C(n26), .ZN(n29) );
  AOI221D0 U90 ( .A1(n35), .A2(search_data[0]), .B1(search_data[13]), .B2(n34), 
        .C(n33), .ZN(n48) );
  AOI221D0 U91 ( .A1(n38), .A2(search_data[14]), .B1(search_data[11]), .B2(n37), .C(n36), .ZN(n47) );
  AOI221D0 U92 ( .A1(n41), .A2(search_data[12]), .B1(search_data[9]), .B2(n40), 
        .C(n39), .ZN(n46) );
  AOI221D0 U93 ( .A1(n44), .A2(search_data[10]), .B1(search_data[25]), .B2(n43), .C(n42), .ZN(n45) );
  AOI221D0 U94 ( .A1(n51), .A2(search_data[7]), .B1(search_data[5]), .B2(n50), 
        .C(n49), .ZN(n65) );
  AOI221D0 U95 ( .A1(n54), .A2(search_data[16]), .B1(search_data[2]), .B2(n53), 
        .C(n52), .ZN(n64) );
  OAI221D0 U96 ( .A1(n57), .A2(search_data[3]), .B1(n56), .B2(search_data[6]), 
        .C(n55), .ZN(n62) );
  OAI221D0 U97 ( .A1(n60), .A2(search_data[1]), .B1(n59), .B2(search_data[4]), 
        .C(n58), .ZN(n61) );
  AO22D0 U98 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U99 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U100 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U101 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U102 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U103 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U104 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U105 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U106 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U107 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U108 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_22 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AN3D0 U4 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results) );
  AO21D0 U5 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  ND4D0 U6 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  NR2D2 U7 ( .A1(reset), .A2(n70), .ZN(n71) );
  CKND2D1 U8 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  AOI21D2 U9 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  OAI22D0 U10 ( .A1(n28), .A2(search_data[18]), .B1(n27), .B2(search_data[15]), 
        .ZN(n26) );
  OAI22D0 U11 ( .A1(n25), .A2(search_data[20]), .B1(n24), .B2(search_data[17]), 
        .ZN(n23) );
  OAI22D0 U12 ( .A1(n38), .A2(search_data[14]), .B1(n37), .B2(search_data[11]), 
        .ZN(n36) );
  OAI22D0 U13 ( .A1(n35), .A2(search_data[0]), .B1(n34), .B2(search_data[13]), 
        .ZN(n33) );
  OAI22D0 U14 ( .A1(n22), .A2(search_data[22]), .B1(n21), .B2(search_data[19]), 
        .ZN(n20) );
  OAI22D0 U15 ( .A1(n41), .A2(search_data[12]), .B1(n40), .B2(search_data[9]), 
        .ZN(n39) );
  OAI22D0 U16 ( .A1(n44), .A2(search_data[10]), .B1(n43), .B2(search_data[25]), 
        .ZN(n42) );
  OAI22D0 U17 ( .A1(n51), .A2(search_data[7]), .B1(n50), .B2(search_data[5]), 
        .ZN(n49) );
  OAI22D0 U18 ( .A1(n54), .A2(search_data[16]), .B1(n53), .B2(search_data[2]), 
        .ZN(n52) );
  AOI22D0 U19 ( .A1(search_data[3]), .A2(n57), .B1(search_data[6]), .B2(n56), 
        .ZN(n55) );
  AOI22D0 U20 ( .A1(search_data[1]), .A2(n60), .B1(search_data[4]), .B2(n59), 
        .ZN(n58) );
  OAI22D0 U21 ( .A1(n3), .A2(search_data[31]), .B1(n2), .B2(search_data[29]), 
        .ZN(n1) );
  OAI22D0 U22 ( .A1(n6), .A2(search_data[30]), .B1(n5), .B2(search_data[27]), 
        .ZN(n4) );
  OAI22D0 U23 ( .A1(n9), .A2(search_data[28]), .B1(n8), .B2(search_data[24]), 
        .ZN(n7) );
  OAI22D0 U24 ( .A1(n12), .A2(search_data[26]), .B1(n11), .B2(search_data[23]), 
        .ZN(n10) );
  OAI22D0 U25 ( .A1(n19), .A2(search_data[8]), .B1(n18), .B2(search_data[21]), 
        .ZN(n17) );
  CKND0 U26 ( .I(read_value[22]), .ZN(n22) );
  CKND0 U27 ( .I(read_value[19]), .ZN(n21) );
  CKND0 U28 ( .I(read_value[23]), .ZN(n11) );
  CKND0 U29 ( .I(read_value[26]), .ZN(n12) );
  CKND0 U30 ( .I(read_value[24]), .ZN(n8) );
  CKND0 U31 ( .I(read_value[8]), .ZN(n19) );
  CKND0 U32 ( .I(read_value[28]), .ZN(n9) );
  CKND0 U33 ( .I(read_value[27]), .ZN(n5) );
  CKND0 U34 ( .I(read_value[30]), .ZN(n6) );
  CKND0 U35 ( .I(read_value[21]), .ZN(n18) );
  CKND0 U36 ( .I(read_value[29]), .ZN(n2) );
  CKND0 U37 ( .I(read_value[31]), .ZN(n3) );
  CKND0 U38 ( .I(read_value[12]), .ZN(n41) );
  CKND0 U39 ( .I(read_value[9]), .ZN(n40) );
  CKND0 U40 ( .I(read_value[10]), .ZN(n44) );
  CKND0 U41 ( .I(read_value[25]), .ZN(n43) );
  CKND0 U42 ( .I(read_value[7]), .ZN(n51) );
  CKND0 U43 ( .I(read_value[5]), .ZN(n50) );
  CKND0 U44 ( .I(read_value[16]), .ZN(n54) );
  CKND0 U45 ( .I(read_value[2]), .ZN(n53) );
  CKND0 U46 ( .I(read_value[3]), .ZN(n57) );
  CKND0 U47 ( .I(read_value[6]), .ZN(n56) );
  CKND0 U48 ( .I(read_value[1]), .ZN(n60) );
  CKND0 U49 ( .I(read_value[4]), .ZN(n59) );
  CKND0 U50 ( .I(read_value[15]), .ZN(n27) );
  CKND0 U51 ( .I(read_value[0]), .ZN(n35) );
  CKND0 U52 ( .I(read_value[18]), .ZN(n28) );
  CKND0 U53 ( .I(read_value[13]), .ZN(n34) );
  CKND0 U54 ( .I(read_value[17]), .ZN(n24) );
  CKND0 U55 ( .I(read_value[14]), .ZN(n38) );
  CKND0 U56 ( .I(read_value[11]), .ZN(n37) );
  CKND0 U57 ( .I(read_value[20]), .ZN(n25) );
  AO22D0 U58 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U59 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U60 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U61 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U62 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U63 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U64 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U65 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), .Z(
        data_i[3]) );
  AO22D0 U66 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U67 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), .Z(
        data_i[2]) );
  AO22D0 U68 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U69 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), .Z(
        data_i[4]) );
  AO22D0 U70 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), .Z(
        data_i[5]) );
  AO22D0 U71 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), .Z(
        data_i[6]) );
  AO22D0 U72 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U73 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U74 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U75 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U76 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U77 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  NR2D1 U78 ( .A1(n62), .A2(n61), .ZN(n63) );
  ND4D1 U79 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .ZN(n67) );
  ND4D1 U80 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .ZN(n68) );
  ND4D1 U81 ( .A1(n16), .A2(n15), .A3(n14), .A4(n13), .ZN(n69) );
  AOI221D0 U82 ( .A1(n3), .A2(search_data[31]), .B1(search_data[29]), .B2(n2), 
        .C(n1), .ZN(n16) );
  AOI221D0 U83 ( .A1(n6), .A2(search_data[30]), .B1(search_data[27]), .B2(n5), 
        .C(n4), .ZN(n15) );
  AOI221D0 U84 ( .A1(n9), .A2(search_data[28]), .B1(search_data[24]), .B2(n8), 
        .C(n7), .ZN(n14) );
  AOI221D0 U85 ( .A1(n12), .A2(search_data[26]), .B1(search_data[23]), .B2(n11), .C(n10), .ZN(n13) );
  AOI221D0 U86 ( .A1(n19), .A2(search_data[8]), .B1(search_data[21]), .B2(n18), 
        .C(n17), .ZN(n32) );
  AOI221D0 U87 ( .A1(n22), .A2(search_data[22]), .B1(search_data[19]), .B2(n21), .C(n20), .ZN(n31) );
  AOI221D0 U88 ( .A1(n25), .A2(search_data[20]), .B1(search_data[17]), .B2(n24), .C(n23), .ZN(n30) );
  AOI221D0 U89 ( .A1(n28), .A2(search_data[18]), .B1(search_data[15]), .B2(n27), .C(n26), .ZN(n29) );
  AOI221D0 U90 ( .A1(n35), .A2(search_data[0]), .B1(search_data[13]), .B2(n34), 
        .C(n33), .ZN(n48) );
  AOI221D0 U91 ( .A1(n38), .A2(search_data[14]), .B1(search_data[11]), .B2(n37), .C(n36), .ZN(n47) );
  AOI221D0 U92 ( .A1(n41), .A2(search_data[12]), .B1(search_data[9]), .B2(n40), 
        .C(n39), .ZN(n46) );
  AOI221D0 U93 ( .A1(n44), .A2(search_data[10]), .B1(search_data[25]), .B2(n43), .C(n42), .ZN(n45) );
  AOI221D0 U94 ( .A1(n51), .A2(search_data[7]), .B1(search_data[5]), .B2(n50), 
        .C(n49), .ZN(n65) );
  AOI221D0 U95 ( .A1(n54), .A2(search_data[16]), .B1(search_data[2]), .B2(n53), 
        .C(n52), .ZN(n64) );
  OAI221D0 U96 ( .A1(n57), .A2(search_data[3]), .B1(n56), .B2(search_data[6]), 
        .C(n55), .ZN(n62) );
  OAI221D0 U97 ( .A1(n60), .A2(search_data[1]), .B1(n59), .B2(search_data[4]), 
        .C(n58), .ZN(n61) );
  AO22D0 U98 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U99 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U100 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U101 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U102 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U103 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U104 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U105 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U106 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U107 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U108 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_23 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AN3D0 U4 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results) );
  ND4D0 U5 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  AO21D0 U6 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U7 ( .A1(reset), .A2(n70), .ZN(n71) );
  CKND2D1 U8 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  AOI21D2 U9 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  OAI22D0 U10 ( .A1(n3), .A2(search_data[31]), .B1(n2), .B2(search_data[29]), 
        .ZN(n1) );
  OAI22D0 U11 ( .A1(n6), .A2(search_data[30]), .B1(n5), .B2(search_data[27]), 
        .ZN(n4) );
  OAI22D0 U12 ( .A1(n9), .A2(search_data[28]), .B1(n8), .B2(search_data[24]), 
        .ZN(n7) );
  OAI22D0 U13 ( .A1(n12), .A2(search_data[26]), .B1(n11), .B2(search_data[23]), 
        .ZN(n10) );
  OAI22D0 U14 ( .A1(n19), .A2(search_data[8]), .B1(n18), .B2(search_data[21]), 
        .ZN(n17) );
  OAI22D0 U15 ( .A1(n22), .A2(search_data[22]), .B1(n21), .B2(search_data[19]), 
        .ZN(n20) );
  OAI22D0 U16 ( .A1(n25), .A2(search_data[20]), .B1(n24), .B2(search_data[17]), 
        .ZN(n23) );
  OAI22D0 U17 ( .A1(n28), .A2(search_data[18]), .B1(n27), .B2(search_data[15]), 
        .ZN(n26) );
  OAI22D0 U18 ( .A1(n35), .A2(search_data[0]), .B1(n34), .B2(search_data[13]), 
        .ZN(n33) );
  OAI22D0 U19 ( .A1(n38), .A2(search_data[14]), .B1(n37), .B2(search_data[11]), 
        .ZN(n36) );
  OAI22D0 U20 ( .A1(n41), .A2(search_data[12]), .B1(n40), .B2(search_data[9]), 
        .ZN(n39) );
  OAI22D0 U21 ( .A1(n44), .A2(search_data[10]), .B1(n43), .B2(search_data[25]), 
        .ZN(n42) );
  OAI22D0 U22 ( .A1(n51), .A2(search_data[7]), .B1(n50), .B2(search_data[5]), 
        .ZN(n49) );
  OAI22D0 U23 ( .A1(n54), .A2(search_data[16]), .B1(n53), .B2(search_data[2]), 
        .ZN(n52) );
  AOI22D0 U24 ( .A1(search_data[3]), .A2(n57), .B1(search_data[6]), .B2(n56), 
        .ZN(n55) );
  AOI22D0 U25 ( .A1(search_data[1]), .A2(n60), .B1(search_data[4]), .B2(n59), 
        .ZN(n58) );
  CKND0 U26 ( .I(read_value[3]), .ZN(n57) );
  CKND0 U27 ( .I(read_value[6]), .ZN(n56) );
  CKND0 U28 ( .I(read_value[1]), .ZN(n60) );
  CKND0 U29 ( .I(read_value[4]), .ZN(n59) );
  CKND0 U30 ( .I(read_value[13]), .ZN(n34) );
  CKND0 U31 ( .I(read_value[0]), .ZN(n35) );
  CKND0 U32 ( .I(read_value[15]), .ZN(n27) );
  CKND0 U33 ( .I(read_value[18]), .ZN(n28) );
  CKND0 U34 ( .I(read_value[17]), .ZN(n24) );
  CKND0 U35 ( .I(read_value[20]), .ZN(n25) );
  CKND0 U36 ( .I(read_value[19]), .ZN(n21) );
  CKND0 U37 ( .I(read_value[22]), .ZN(n22) );
  CKND0 U38 ( .I(read_value[21]), .ZN(n18) );
  CKND0 U39 ( .I(read_value[8]), .ZN(n19) );
  CKND0 U40 ( .I(read_value[23]), .ZN(n11) );
  CKND0 U41 ( .I(read_value[26]), .ZN(n12) );
  CKND0 U42 ( .I(read_value[24]), .ZN(n8) );
  CKND0 U43 ( .I(read_value[28]), .ZN(n9) );
  CKND0 U44 ( .I(read_value[27]), .ZN(n5) );
  CKND0 U45 ( .I(read_value[30]), .ZN(n6) );
  CKND0 U46 ( .I(read_value[29]), .ZN(n2) );
  CKND0 U47 ( .I(read_value[31]), .ZN(n3) );
  CKND0 U48 ( .I(read_value[25]), .ZN(n43) );
  CKND0 U49 ( .I(read_value[10]), .ZN(n44) );
  CKND0 U50 ( .I(read_value[5]), .ZN(n50) );
  CKND0 U51 ( .I(read_value[9]), .ZN(n40) );
  CKND0 U52 ( .I(read_value[12]), .ZN(n41) );
  CKND0 U53 ( .I(read_value[7]), .ZN(n51) );
  CKND0 U54 ( .I(read_value[14]), .ZN(n38) );
  CKND0 U55 ( .I(read_value[2]), .ZN(n53) );
  CKND0 U56 ( .I(read_value[16]), .ZN(n54) );
  CKND0 U57 ( .I(read_value[11]), .ZN(n37) );
  AO22D0 U58 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U59 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U60 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U61 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U62 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U63 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U64 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U65 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U66 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U67 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U68 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U69 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), .Z(
        data_i[2]) );
  AO22D0 U70 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U71 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), .Z(
        data_i[6]) );
  AO22D0 U72 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), .Z(
        data_i[5]) );
  AO22D0 U73 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), .Z(
        data_i[4]) );
  AO22D0 U74 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), .Z(
        data_i[3]) );
  AO22D0 U75 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U76 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U77 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  NR2D1 U78 ( .A1(n62), .A2(n61), .ZN(n63) );
  ND4D1 U79 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .ZN(n67) );
  ND4D1 U80 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .ZN(n68) );
  ND4D1 U81 ( .A1(n16), .A2(n15), .A3(n14), .A4(n13), .ZN(n69) );
  AOI221D0 U82 ( .A1(n3), .A2(search_data[31]), .B1(search_data[29]), .B2(n2), 
        .C(n1), .ZN(n16) );
  AOI221D0 U83 ( .A1(n6), .A2(search_data[30]), .B1(search_data[27]), .B2(n5), 
        .C(n4), .ZN(n15) );
  AOI221D0 U84 ( .A1(n9), .A2(search_data[28]), .B1(search_data[24]), .B2(n8), 
        .C(n7), .ZN(n14) );
  AOI221D0 U85 ( .A1(n12), .A2(search_data[26]), .B1(search_data[23]), .B2(n11), .C(n10), .ZN(n13) );
  AOI221D0 U86 ( .A1(n19), .A2(search_data[8]), .B1(search_data[21]), .B2(n18), 
        .C(n17), .ZN(n32) );
  AOI221D0 U87 ( .A1(n22), .A2(search_data[22]), .B1(search_data[19]), .B2(n21), .C(n20), .ZN(n31) );
  AOI221D0 U88 ( .A1(n25), .A2(search_data[20]), .B1(search_data[17]), .B2(n24), .C(n23), .ZN(n30) );
  AOI221D0 U89 ( .A1(n28), .A2(search_data[18]), .B1(search_data[15]), .B2(n27), .C(n26), .ZN(n29) );
  AOI221D0 U90 ( .A1(n35), .A2(search_data[0]), .B1(search_data[13]), .B2(n34), 
        .C(n33), .ZN(n48) );
  AOI221D0 U91 ( .A1(n38), .A2(search_data[14]), .B1(search_data[11]), .B2(n37), .C(n36), .ZN(n47) );
  AOI221D0 U92 ( .A1(n41), .A2(search_data[12]), .B1(search_data[9]), .B2(n40), 
        .C(n39), .ZN(n46) );
  AOI221D0 U93 ( .A1(n44), .A2(search_data[10]), .B1(search_data[25]), .B2(n43), .C(n42), .ZN(n45) );
  AOI221D0 U94 ( .A1(n51), .A2(search_data[7]), .B1(search_data[5]), .B2(n50), 
        .C(n49), .ZN(n65) );
  AOI221D0 U95 ( .A1(n54), .A2(search_data[16]), .B1(search_data[2]), .B2(n53), 
        .C(n52), .ZN(n64) );
  OAI221D0 U96 ( .A1(n57), .A2(search_data[3]), .B1(n56), .B2(search_data[6]), 
        .C(n55), .ZN(n62) );
  OAI221D0 U97 ( .A1(n60), .A2(search_data[1]), .B1(n59), .B2(search_data[4]), 
        .C(n58), .ZN(n61) );
  AO22D0 U98 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U99 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U100 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U101 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U102 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U103 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U104 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U105 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U106 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U107 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U108 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_24 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AN3D0 U4 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results) );
  ND4D0 U5 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  AO21D0 U6 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U7 ( .A1(reset), .A2(n70), .ZN(n71) );
  CKND2D1 U8 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  AOI21D2 U9 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  AOI22D0 U10 ( .A1(search_data[1]), .A2(n60), .B1(search_data[4]), .B2(n59), 
        .ZN(n58) );
  AOI22D0 U11 ( .A1(search_data[3]), .A2(n57), .B1(search_data[6]), .B2(n56), 
        .ZN(n55) );
  OAI22D0 U12 ( .A1(n54), .A2(search_data[16]), .B1(n53), .B2(search_data[2]), 
        .ZN(n52) );
  OAI22D0 U13 ( .A1(n51), .A2(search_data[7]), .B1(n50), .B2(search_data[5]), 
        .ZN(n49) );
  OAI22D0 U14 ( .A1(n44), .A2(search_data[10]), .B1(n43), .B2(search_data[25]), 
        .ZN(n42) );
  OAI22D0 U15 ( .A1(n41), .A2(search_data[12]), .B1(n40), .B2(search_data[9]), 
        .ZN(n39) );
  OAI22D0 U16 ( .A1(n38), .A2(search_data[14]), .B1(n37), .B2(search_data[11]), 
        .ZN(n36) );
  OAI22D0 U17 ( .A1(n3), .A2(search_data[31]), .B1(n2), .B2(search_data[29]), 
        .ZN(n1) );
  OAI22D0 U18 ( .A1(n35), .A2(search_data[0]), .B1(n34), .B2(search_data[13]), 
        .ZN(n33) );
  OAI22D0 U19 ( .A1(n6), .A2(search_data[30]), .B1(n5), .B2(search_data[27]), 
        .ZN(n4) );
  OAI22D0 U20 ( .A1(n28), .A2(search_data[18]), .B1(n27), .B2(search_data[15]), 
        .ZN(n26) );
  OAI22D0 U21 ( .A1(n9), .A2(search_data[28]), .B1(n8), .B2(search_data[24]), 
        .ZN(n7) );
  OAI22D0 U22 ( .A1(n25), .A2(search_data[20]), .B1(n24), .B2(search_data[17]), 
        .ZN(n23) );
  OAI22D0 U23 ( .A1(n22), .A2(search_data[22]), .B1(n21), .B2(search_data[19]), 
        .ZN(n20) );
  OAI22D0 U24 ( .A1(n12), .A2(search_data[26]), .B1(n11), .B2(search_data[23]), 
        .ZN(n10) );
  OAI22D0 U25 ( .A1(n19), .A2(search_data[8]), .B1(n18), .B2(search_data[21]), 
        .ZN(n17) );
  CKND0 U26 ( .I(read_value[4]), .ZN(n59) );
  CKND0 U27 ( .I(read_value[1]), .ZN(n60) );
  CKND0 U28 ( .I(read_value[6]), .ZN(n56) );
  CKND0 U29 ( .I(read_value[3]), .ZN(n57) );
  CKND0 U30 ( .I(read_value[2]), .ZN(n53) );
  CKND0 U31 ( .I(read_value[16]), .ZN(n54) );
  CKND0 U32 ( .I(read_value[5]), .ZN(n50) );
  CKND0 U33 ( .I(read_value[7]), .ZN(n51) );
  CKND0 U34 ( .I(read_value[25]), .ZN(n43) );
  CKND0 U35 ( .I(read_value[10]), .ZN(n44) );
  CKND0 U36 ( .I(read_value[9]), .ZN(n40) );
  CKND0 U37 ( .I(read_value[12]), .ZN(n41) );
  CKND0 U38 ( .I(read_value[11]), .ZN(n37) );
  CKND0 U39 ( .I(read_value[14]), .ZN(n38) );
  CKND0 U40 ( .I(read_value[31]), .ZN(n3) );
  CKND0 U41 ( .I(read_value[13]), .ZN(n34) );
  CKND0 U42 ( .I(read_value[29]), .ZN(n2) );
  CKND0 U43 ( .I(read_value[0]), .ZN(n35) );
  CKND0 U44 ( .I(read_value[30]), .ZN(n6) );
  CKND0 U45 ( .I(read_value[15]), .ZN(n27) );
  CKND0 U46 ( .I(read_value[18]), .ZN(n28) );
  CKND0 U47 ( .I(read_value[27]), .ZN(n5) );
  CKND0 U48 ( .I(read_value[17]), .ZN(n24) );
  CKND0 U49 ( .I(read_value[20]), .ZN(n25) );
  CKND0 U50 ( .I(read_value[28]), .ZN(n9) );
  CKND0 U51 ( .I(read_value[24]), .ZN(n8) );
  CKND0 U52 ( .I(read_value[19]), .ZN(n21) );
  CKND0 U53 ( .I(read_value[22]), .ZN(n22) );
  CKND0 U54 ( .I(read_value[26]), .ZN(n12) );
  CKND0 U55 ( .I(read_value[21]), .ZN(n18) );
  CKND0 U56 ( .I(read_value[8]), .ZN(n19) );
  CKND0 U57 ( .I(read_value[23]), .ZN(n11) );
  AO22D0 U58 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), .Z(
        data_i[5]) );
  AO22D0 U59 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U60 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), .Z(
        data_i[4]) );
  AO22D0 U61 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U62 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U63 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), .Z(
        data_i[2]) );
  AO22D0 U64 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U65 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), .Z(
        data_i[6]) );
  AO22D0 U66 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U67 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U68 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U69 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U70 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U71 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U72 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U73 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), .Z(
        data_i[3]) );
  AO22D0 U74 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U75 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U76 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U77 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  NR2D1 U78 ( .A1(n62), .A2(n61), .ZN(n63) );
  ND4D1 U79 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .ZN(n67) );
  ND4D1 U80 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .ZN(n68) );
  ND4D1 U81 ( .A1(n16), .A2(n15), .A3(n14), .A4(n13), .ZN(n69) );
  AOI221D0 U82 ( .A1(n3), .A2(search_data[31]), .B1(search_data[29]), .B2(n2), 
        .C(n1), .ZN(n16) );
  AOI221D0 U83 ( .A1(n6), .A2(search_data[30]), .B1(search_data[27]), .B2(n5), 
        .C(n4), .ZN(n15) );
  AOI221D0 U84 ( .A1(n9), .A2(search_data[28]), .B1(search_data[24]), .B2(n8), 
        .C(n7), .ZN(n14) );
  AOI221D0 U85 ( .A1(n12), .A2(search_data[26]), .B1(search_data[23]), .B2(n11), .C(n10), .ZN(n13) );
  AOI221D0 U86 ( .A1(n19), .A2(search_data[8]), .B1(search_data[21]), .B2(n18), 
        .C(n17), .ZN(n32) );
  AOI221D0 U87 ( .A1(n22), .A2(search_data[22]), .B1(search_data[19]), .B2(n21), .C(n20), .ZN(n31) );
  AOI221D0 U88 ( .A1(n25), .A2(search_data[20]), .B1(search_data[17]), .B2(n24), .C(n23), .ZN(n30) );
  AOI221D0 U89 ( .A1(n28), .A2(search_data[18]), .B1(search_data[15]), .B2(n27), .C(n26), .ZN(n29) );
  AOI221D0 U90 ( .A1(n35), .A2(search_data[0]), .B1(search_data[13]), .B2(n34), 
        .C(n33), .ZN(n48) );
  AOI221D0 U91 ( .A1(n38), .A2(search_data[14]), .B1(search_data[11]), .B2(n37), .C(n36), .ZN(n47) );
  AOI221D0 U92 ( .A1(n41), .A2(search_data[12]), .B1(search_data[9]), .B2(n40), 
        .C(n39), .ZN(n46) );
  AOI221D0 U93 ( .A1(n44), .A2(search_data[10]), .B1(search_data[25]), .B2(n43), .C(n42), .ZN(n45) );
  AOI221D0 U94 ( .A1(n51), .A2(search_data[7]), .B1(search_data[5]), .B2(n50), 
        .C(n49), .ZN(n65) );
  AOI221D0 U95 ( .A1(n54), .A2(search_data[16]), .B1(search_data[2]), .B2(n53), 
        .C(n52), .ZN(n64) );
  OAI221D0 U96 ( .A1(n57), .A2(search_data[3]), .B1(n56), .B2(search_data[6]), 
        .C(n55), .ZN(n62) );
  OAI221D0 U97 ( .A1(n60), .A2(search_data[1]), .B1(n59), .B2(search_data[4]), 
        .C(n58), .ZN(n61) );
  AO22D0 U98 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U99 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U100 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U101 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U102 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U103 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U104 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U105 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U106 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U107 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U108 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_25 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AN3D0 U4 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results) );
  ND4D0 U5 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  AO21D0 U6 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U7 ( .A1(reset), .A2(n70), .ZN(n71) );
  CKND2D1 U8 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  AOI21D2 U9 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  AOI22D0 U10 ( .A1(search_data[1]), .A2(n60), .B1(search_data[4]), .B2(n59), 
        .ZN(n58) );
  AOI22D0 U11 ( .A1(search_data[3]), .A2(n57), .B1(search_data[6]), .B2(n56), 
        .ZN(n55) );
  OAI22D0 U12 ( .A1(n54), .A2(search_data[16]), .B1(n53), .B2(search_data[2]), 
        .ZN(n52) );
  OAI22D0 U13 ( .A1(n51), .A2(search_data[7]), .B1(n50), .B2(search_data[5]), 
        .ZN(n49) );
  OAI22D0 U14 ( .A1(n44), .A2(search_data[10]), .B1(n43), .B2(search_data[25]), 
        .ZN(n42) );
  OAI22D0 U15 ( .A1(n41), .A2(search_data[12]), .B1(n40), .B2(search_data[9]), 
        .ZN(n39) );
  OAI22D0 U16 ( .A1(n38), .A2(search_data[14]), .B1(n37), .B2(search_data[11]), 
        .ZN(n36) );
  OAI22D0 U17 ( .A1(n35), .A2(search_data[0]), .B1(n34), .B2(search_data[13]), 
        .ZN(n33) );
  OAI22D0 U18 ( .A1(n28), .A2(search_data[18]), .B1(n27), .B2(search_data[15]), 
        .ZN(n26) );
  OAI22D0 U19 ( .A1(n25), .A2(search_data[20]), .B1(n24), .B2(search_data[17]), 
        .ZN(n23) );
  OAI22D0 U20 ( .A1(n22), .A2(search_data[22]), .B1(n21), .B2(search_data[19]), 
        .ZN(n20) );
  OAI22D0 U21 ( .A1(n19), .A2(search_data[8]), .B1(n18), .B2(search_data[21]), 
        .ZN(n17) );
  OAI22D0 U22 ( .A1(n12), .A2(search_data[26]), .B1(n11), .B2(search_data[23]), 
        .ZN(n10) );
  OAI22D0 U23 ( .A1(n9), .A2(search_data[28]), .B1(n8), .B2(search_data[24]), 
        .ZN(n7) );
  OAI22D0 U24 ( .A1(n6), .A2(search_data[30]), .B1(n5), .B2(search_data[27]), 
        .ZN(n4) );
  OAI22D0 U25 ( .A1(n3), .A2(search_data[31]), .B1(n2), .B2(search_data[29]), 
        .ZN(n1) );
  CKND0 U26 ( .I(read_value[4]), .ZN(n59) );
  CKND0 U27 ( .I(read_value[1]), .ZN(n60) );
  CKND0 U28 ( .I(read_value[6]), .ZN(n56) );
  CKND0 U29 ( .I(read_value[3]), .ZN(n57) );
  CKND0 U30 ( .I(read_value[29]), .ZN(n2) );
  CKND0 U31 ( .I(read_value[31]), .ZN(n3) );
  CKND0 U32 ( .I(read_value[2]), .ZN(n53) );
  CKND0 U33 ( .I(read_value[16]), .ZN(n54) );
  CKND0 U34 ( .I(read_value[5]), .ZN(n50) );
  CKND0 U35 ( .I(read_value[7]), .ZN(n51) );
  CKND0 U36 ( .I(read_value[25]), .ZN(n43) );
  CKND0 U37 ( .I(read_value[10]), .ZN(n44) );
  CKND0 U38 ( .I(read_value[9]), .ZN(n40) );
  CKND0 U39 ( .I(read_value[12]), .ZN(n41) );
  CKND0 U40 ( .I(read_value[11]), .ZN(n37) );
  CKND0 U41 ( .I(read_value[14]), .ZN(n38) );
  CKND0 U42 ( .I(read_value[13]), .ZN(n34) );
  CKND0 U43 ( .I(read_value[0]), .ZN(n35) );
  CKND0 U44 ( .I(read_value[15]), .ZN(n27) );
  CKND0 U45 ( .I(read_value[18]), .ZN(n28) );
  CKND0 U46 ( .I(read_value[17]), .ZN(n24) );
  CKND0 U47 ( .I(read_value[20]), .ZN(n25) );
  CKND0 U48 ( .I(read_value[19]), .ZN(n21) );
  CKND0 U49 ( .I(read_value[22]), .ZN(n22) );
  CKND0 U50 ( .I(read_value[21]), .ZN(n18) );
  CKND0 U51 ( .I(read_value[8]), .ZN(n19) );
  CKND0 U52 ( .I(read_value[23]), .ZN(n11) );
  CKND0 U53 ( .I(read_value[26]), .ZN(n12) );
  CKND0 U54 ( .I(read_value[24]), .ZN(n8) );
  CKND0 U55 ( .I(read_value[28]), .ZN(n9) );
  CKND0 U56 ( .I(read_value[27]), .ZN(n5) );
  CKND0 U57 ( .I(read_value[30]), .ZN(n6) );
  AO22D0 U58 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U59 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U60 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U61 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), .Z(
        data_i[2]) );
  AO22D0 U62 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), .Z(
        data_i[3]) );
  AO22D0 U63 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), .Z(
        data_i[4]) );
  AO22D0 U64 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), .Z(
        data_i[5]) );
  AO22D0 U65 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), .Z(
        data_i[6]) );
  AO22D0 U66 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U67 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U68 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U69 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U70 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U71 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U72 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U73 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U74 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U75 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U76 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U77 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  NR2D1 U78 ( .A1(n62), .A2(n61), .ZN(n63) );
  ND4D1 U79 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .ZN(n67) );
  ND4D1 U80 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .ZN(n68) );
  ND4D1 U81 ( .A1(n16), .A2(n15), .A3(n14), .A4(n13), .ZN(n69) );
  AOI221D0 U82 ( .A1(n3), .A2(search_data[31]), .B1(search_data[29]), .B2(n2), 
        .C(n1), .ZN(n16) );
  AOI221D0 U83 ( .A1(n6), .A2(search_data[30]), .B1(search_data[27]), .B2(n5), 
        .C(n4), .ZN(n15) );
  AOI221D0 U84 ( .A1(n9), .A2(search_data[28]), .B1(search_data[24]), .B2(n8), 
        .C(n7), .ZN(n14) );
  AOI221D0 U85 ( .A1(n12), .A2(search_data[26]), .B1(search_data[23]), .B2(n11), .C(n10), .ZN(n13) );
  AOI221D0 U86 ( .A1(n19), .A2(search_data[8]), .B1(search_data[21]), .B2(n18), 
        .C(n17), .ZN(n32) );
  AOI221D0 U87 ( .A1(n22), .A2(search_data[22]), .B1(search_data[19]), .B2(n21), .C(n20), .ZN(n31) );
  AOI221D0 U88 ( .A1(n25), .A2(search_data[20]), .B1(search_data[17]), .B2(n24), .C(n23), .ZN(n30) );
  AOI221D0 U89 ( .A1(n28), .A2(search_data[18]), .B1(search_data[15]), .B2(n27), .C(n26), .ZN(n29) );
  AOI221D0 U90 ( .A1(n35), .A2(search_data[0]), .B1(search_data[13]), .B2(n34), 
        .C(n33), .ZN(n48) );
  AOI221D0 U91 ( .A1(n38), .A2(search_data[14]), .B1(search_data[11]), .B2(n37), .C(n36), .ZN(n47) );
  AOI221D0 U92 ( .A1(n41), .A2(search_data[12]), .B1(search_data[9]), .B2(n40), 
        .C(n39), .ZN(n46) );
  AOI221D0 U93 ( .A1(n44), .A2(search_data[10]), .B1(search_data[25]), .B2(n43), .C(n42), .ZN(n45) );
  AOI221D0 U94 ( .A1(n51), .A2(search_data[7]), .B1(search_data[5]), .B2(n50), 
        .C(n49), .ZN(n65) );
  AOI221D0 U95 ( .A1(n54), .A2(search_data[16]), .B1(search_data[2]), .B2(n53), 
        .C(n52), .ZN(n64) );
  OAI221D0 U96 ( .A1(n57), .A2(search_data[3]), .B1(n56), .B2(search_data[6]), 
        .C(n55), .ZN(n62) );
  OAI221D0 U97 ( .A1(n60), .A2(search_data[1]), .B1(n59), .B2(search_data[4]), 
        .C(n58), .ZN(n61) );
  AO22D0 U98 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U99 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U100 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U101 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U102 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U103 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U104 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U105 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U106 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U107 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U108 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_26 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AN3D0 U4 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results) );
  AO21D0 U5 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  ND4D0 U6 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  NR2D2 U7 ( .A1(reset), .A2(n70), .ZN(n71) );
  CKND2D1 U8 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  AOI21D2 U9 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  OAI22D0 U10 ( .A1(n51), .A2(search_data[7]), .B1(n50), .B2(search_data[5]), 
        .ZN(n49) );
  OAI22D0 U11 ( .A1(n54), .A2(search_data[16]), .B1(n53), .B2(search_data[2]), 
        .ZN(n52) );
  AOI22D0 U12 ( .A1(search_data[3]), .A2(n57), .B1(search_data[6]), .B2(n56), 
        .ZN(n55) );
  AOI22D0 U13 ( .A1(search_data[1]), .A2(n60), .B1(search_data[4]), .B2(n59), 
        .ZN(n58) );
  OAI22D0 U14 ( .A1(n44), .A2(search_data[10]), .B1(n43), .B2(search_data[25]), 
        .ZN(n42) );
  OAI22D0 U15 ( .A1(n3), .A2(search_data[31]), .B1(n2), .B2(search_data[29]), 
        .ZN(n1) );
  OAI22D0 U16 ( .A1(n6), .A2(search_data[30]), .B1(n5), .B2(search_data[27]), 
        .ZN(n4) );
  OAI22D0 U17 ( .A1(n9), .A2(search_data[28]), .B1(n8), .B2(search_data[24]), 
        .ZN(n7) );
  OAI22D0 U18 ( .A1(n12), .A2(search_data[26]), .B1(n11), .B2(search_data[23]), 
        .ZN(n10) );
  OAI22D0 U19 ( .A1(n19), .A2(search_data[8]), .B1(n18), .B2(search_data[21]), 
        .ZN(n17) );
  OAI22D0 U20 ( .A1(n22), .A2(search_data[22]), .B1(n21), .B2(search_data[19]), 
        .ZN(n20) );
  OAI22D0 U21 ( .A1(n25), .A2(search_data[20]), .B1(n24), .B2(search_data[17]), 
        .ZN(n23) );
  OAI22D0 U22 ( .A1(n28), .A2(search_data[18]), .B1(n27), .B2(search_data[15]), 
        .ZN(n26) );
  OAI22D0 U23 ( .A1(n35), .A2(search_data[0]), .B1(n34), .B2(search_data[13]), 
        .ZN(n33) );
  OAI22D0 U24 ( .A1(n38), .A2(search_data[14]), .B1(n37), .B2(search_data[11]), 
        .ZN(n36) );
  OAI22D0 U25 ( .A1(n41), .A2(search_data[12]), .B1(n40), .B2(search_data[9]), 
        .ZN(n39) );
  CKND0 U26 ( .I(read_value[15]), .ZN(n27) );
  CKND0 U27 ( .I(read_value[0]), .ZN(n35) );
  CKND0 U28 ( .I(read_value[13]), .ZN(n34) );
  CKND0 U29 ( .I(read_value[14]), .ZN(n38) );
  CKND0 U30 ( .I(read_value[11]), .ZN(n37) );
  CKND0 U31 ( .I(read_value[12]), .ZN(n41) );
  CKND0 U32 ( .I(read_value[9]), .ZN(n40) );
  CKND0 U33 ( .I(read_value[10]), .ZN(n44) );
  CKND0 U34 ( .I(read_value[25]), .ZN(n43) );
  CKND0 U35 ( .I(read_value[7]), .ZN(n51) );
  CKND0 U36 ( .I(read_value[5]), .ZN(n50) );
  CKND0 U37 ( .I(read_value[16]), .ZN(n54) );
  CKND0 U38 ( .I(read_value[2]), .ZN(n53) );
  CKND0 U39 ( .I(read_value[3]), .ZN(n57) );
  CKND0 U40 ( .I(read_value[6]), .ZN(n56) );
  CKND0 U41 ( .I(read_value[1]), .ZN(n60) );
  CKND0 U42 ( .I(read_value[4]), .ZN(n59) );
  CKND0 U43 ( .I(read_value[18]), .ZN(n28) );
  CKND0 U44 ( .I(read_value[31]), .ZN(n3) );
  CKND0 U45 ( .I(read_value[29]), .ZN(n2) );
  CKND0 U46 ( .I(read_value[30]), .ZN(n6) );
  CKND0 U47 ( .I(read_value[27]), .ZN(n5) );
  CKND0 U48 ( .I(read_value[28]), .ZN(n9) );
  CKND0 U49 ( .I(read_value[24]), .ZN(n8) );
  CKND0 U50 ( .I(read_value[26]), .ZN(n12) );
  CKND0 U51 ( .I(read_value[23]), .ZN(n11) );
  CKND0 U52 ( .I(read_value[8]), .ZN(n19) );
  CKND0 U53 ( .I(read_value[21]), .ZN(n18) );
  CKND0 U54 ( .I(read_value[22]), .ZN(n22) );
  CKND0 U55 ( .I(read_value[19]), .ZN(n21) );
  CKND0 U56 ( .I(read_value[20]), .ZN(n25) );
  CKND0 U57 ( .I(read_value[17]), .ZN(n24) );
  AO22D0 U58 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U59 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U60 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U61 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U62 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U63 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U64 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U65 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U66 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U67 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U68 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U69 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U70 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U71 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), .Z(
        data_i[6]) );
  AO22D0 U72 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), .Z(
        data_i[5]) );
  AO22D0 U73 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), .Z(
        data_i[4]) );
  AO22D0 U74 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), .Z(
        data_i[3]) );
  AO22D0 U75 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), .Z(
        data_i[2]) );
  AO22D0 U76 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U77 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  NR2D1 U78 ( .A1(n62), .A2(n61), .ZN(n63) );
  ND4D1 U79 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .ZN(n67) );
  ND4D1 U80 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .ZN(n68) );
  ND4D1 U81 ( .A1(n16), .A2(n15), .A3(n14), .A4(n13), .ZN(n69) );
  AOI221D0 U82 ( .A1(n3), .A2(search_data[31]), .B1(search_data[29]), .B2(n2), 
        .C(n1), .ZN(n16) );
  AOI221D0 U83 ( .A1(n6), .A2(search_data[30]), .B1(search_data[27]), .B2(n5), 
        .C(n4), .ZN(n15) );
  AOI221D0 U84 ( .A1(n9), .A2(search_data[28]), .B1(search_data[24]), .B2(n8), 
        .C(n7), .ZN(n14) );
  AOI221D0 U85 ( .A1(n12), .A2(search_data[26]), .B1(search_data[23]), .B2(n11), .C(n10), .ZN(n13) );
  AOI221D0 U86 ( .A1(n19), .A2(search_data[8]), .B1(search_data[21]), .B2(n18), 
        .C(n17), .ZN(n32) );
  AOI221D0 U87 ( .A1(n22), .A2(search_data[22]), .B1(search_data[19]), .B2(n21), .C(n20), .ZN(n31) );
  AOI221D0 U88 ( .A1(n25), .A2(search_data[20]), .B1(search_data[17]), .B2(n24), .C(n23), .ZN(n30) );
  AOI221D0 U89 ( .A1(n28), .A2(search_data[18]), .B1(search_data[15]), .B2(n27), .C(n26), .ZN(n29) );
  AOI221D0 U90 ( .A1(n35), .A2(search_data[0]), .B1(search_data[13]), .B2(n34), 
        .C(n33), .ZN(n48) );
  AOI221D0 U91 ( .A1(n38), .A2(search_data[14]), .B1(search_data[11]), .B2(n37), .C(n36), .ZN(n47) );
  AOI221D0 U92 ( .A1(n41), .A2(search_data[12]), .B1(search_data[9]), .B2(n40), 
        .C(n39), .ZN(n46) );
  AOI221D0 U93 ( .A1(n44), .A2(search_data[10]), .B1(search_data[25]), .B2(n43), .C(n42), .ZN(n45) );
  AOI221D0 U94 ( .A1(n51), .A2(search_data[7]), .B1(search_data[5]), .B2(n50), 
        .C(n49), .ZN(n65) );
  AOI221D0 U95 ( .A1(n54), .A2(search_data[16]), .B1(search_data[2]), .B2(n53), 
        .C(n52), .ZN(n64) );
  OAI221D0 U96 ( .A1(n57), .A2(search_data[3]), .B1(n56), .B2(search_data[6]), 
        .C(n55), .ZN(n62) );
  OAI221D0 U97 ( .A1(n60), .A2(search_data[1]), .B1(n59), .B2(search_data[4]), 
        .C(n58), .ZN(n61) );
  AO22D0 U98 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U99 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U100 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U101 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U102 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U103 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U104 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U105 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U106 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U107 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U108 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_27 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AN3D0 U4 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results) );
  ND4D0 U5 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  AO21D0 U6 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U7 ( .A1(reset), .A2(n70), .ZN(n71) );
  CKND2D1 U8 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  AOI21D2 U9 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  OAI22D0 U10 ( .A1(n3), .A2(search_data[31]), .B1(n2), .B2(search_data[29]), 
        .ZN(n1) );
  OAI22D0 U11 ( .A1(n6), .A2(search_data[30]), .B1(n5), .B2(search_data[27]), 
        .ZN(n4) );
  OAI22D0 U12 ( .A1(n9), .A2(search_data[28]), .B1(n8), .B2(search_data[24]), 
        .ZN(n7) );
  OAI22D0 U13 ( .A1(n12), .A2(search_data[26]), .B1(n11), .B2(search_data[23]), 
        .ZN(n10) );
  OAI22D0 U14 ( .A1(n19), .A2(search_data[8]), .B1(n18), .B2(search_data[21]), 
        .ZN(n17) );
  OAI22D0 U15 ( .A1(n22), .A2(search_data[22]), .B1(n21), .B2(search_data[19]), 
        .ZN(n20) );
  OAI22D0 U16 ( .A1(n25), .A2(search_data[20]), .B1(n24), .B2(search_data[17]), 
        .ZN(n23) );
  OAI22D0 U17 ( .A1(n28), .A2(search_data[18]), .B1(n27), .B2(search_data[15]), 
        .ZN(n26) );
  OAI22D0 U18 ( .A1(n35), .A2(search_data[0]), .B1(n34), .B2(search_data[13]), 
        .ZN(n33) );
  OAI22D0 U19 ( .A1(n38), .A2(search_data[14]), .B1(n37), .B2(search_data[11]), 
        .ZN(n36) );
  OAI22D0 U20 ( .A1(n41), .A2(search_data[12]), .B1(n40), .B2(search_data[9]), 
        .ZN(n39) );
  OAI22D0 U21 ( .A1(n44), .A2(search_data[10]), .B1(n43), .B2(search_data[25]), 
        .ZN(n42) );
  OAI22D0 U22 ( .A1(n51), .A2(search_data[7]), .B1(n50), .B2(search_data[5]), 
        .ZN(n49) );
  OAI22D0 U23 ( .A1(n54), .A2(search_data[16]), .B1(n53), .B2(search_data[2]), 
        .ZN(n52) );
  AOI22D0 U24 ( .A1(search_data[3]), .A2(n57), .B1(search_data[6]), .B2(n56), 
        .ZN(n55) );
  AOI22D0 U25 ( .A1(search_data[1]), .A2(n60), .B1(search_data[4]), .B2(n59), 
        .ZN(n58) );
  CKND0 U26 ( .I(read_value[31]), .ZN(n3) );
  CKND0 U27 ( .I(read_value[29]), .ZN(n2) );
  CKND0 U28 ( .I(read_value[9]), .ZN(n40) );
  CKND0 U29 ( .I(read_value[10]), .ZN(n44) );
  CKND0 U30 ( .I(read_value[25]), .ZN(n43) );
  CKND0 U31 ( .I(read_value[7]), .ZN(n51) );
  CKND0 U32 ( .I(read_value[5]), .ZN(n50) );
  CKND0 U33 ( .I(read_value[16]), .ZN(n54) );
  CKND0 U34 ( .I(read_value[2]), .ZN(n53) );
  CKND0 U35 ( .I(read_value[3]), .ZN(n57) );
  CKND0 U36 ( .I(read_value[6]), .ZN(n56) );
  CKND0 U37 ( .I(read_value[12]), .ZN(n41) );
  CKND0 U38 ( .I(read_value[1]), .ZN(n60) );
  CKND0 U39 ( .I(read_value[4]), .ZN(n59) );
  CKND0 U40 ( .I(read_value[30]), .ZN(n6) );
  CKND0 U41 ( .I(read_value[27]), .ZN(n5) );
  CKND0 U42 ( .I(read_value[28]), .ZN(n9) );
  CKND0 U43 ( .I(read_value[24]), .ZN(n8) );
  CKND0 U44 ( .I(read_value[26]), .ZN(n12) );
  CKND0 U45 ( .I(read_value[23]), .ZN(n11) );
  CKND0 U46 ( .I(read_value[8]), .ZN(n19) );
  CKND0 U47 ( .I(read_value[21]), .ZN(n18) );
  CKND0 U48 ( .I(read_value[22]), .ZN(n22) );
  CKND0 U49 ( .I(read_value[19]), .ZN(n21) );
  CKND0 U50 ( .I(read_value[20]), .ZN(n25) );
  CKND0 U51 ( .I(read_value[17]), .ZN(n24) );
  CKND0 U52 ( .I(read_value[18]), .ZN(n28) );
  CKND0 U53 ( .I(read_value[15]), .ZN(n27) );
  CKND0 U54 ( .I(read_value[0]), .ZN(n35) );
  CKND0 U55 ( .I(read_value[13]), .ZN(n34) );
  CKND0 U56 ( .I(read_value[14]), .ZN(n38) );
  CKND0 U57 ( .I(read_value[11]), .ZN(n37) );
  AO22D0 U58 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U59 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U60 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U61 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U62 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U63 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U64 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U65 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U66 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U67 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U68 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U69 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U70 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U71 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), .Z(
        data_i[6]) );
  AO22D0 U72 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), .Z(
        data_i[5]) );
  AO22D0 U73 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), .Z(
        data_i[4]) );
  AO22D0 U74 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), .Z(
        data_i[3]) );
  AO22D0 U75 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), .Z(
        data_i[2]) );
  AO22D0 U76 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U77 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  NR2D1 U78 ( .A1(n62), .A2(n61), .ZN(n63) );
  ND4D1 U79 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .ZN(n67) );
  ND4D1 U80 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .ZN(n68) );
  ND4D1 U81 ( .A1(n16), .A2(n15), .A3(n14), .A4(n13), .ZN(n69) );
  AOI221D0 U82 ( .A1(n3), .A2(search_data[31]), .B1(search_data[29]), .B2(n2), 
        .C(n1), .ZN(n16) );
  AOI221D0 U83 ( .A1(n6), .A2(search_data[30]), .B1(search_data[27]), .B2(n5), 
        .C(n4), .ZN(n15) );
  AOI221D0 U84 ( .A1(n9), .A2(search_data[28]), .B1(search_data[24]), .B2(n8), 
        .C(n7), .ZN(n14) );
  AOI221D0 U85 ( .A1(n12), .A2(search_data[26]), .B1(search_data[23]), .B2(n11), .C(n10), .ZN(n13) );
  AOI221D0 U86 ( .A1(n19), .A2(search_data[8]), .B1(search_data[21]), .B2(n18), 
        .C(n17), .ZN(n32) );
  AOI221D0 U87 ( .A1(n22), .A2(search_data[22]), .B1(search_data[19]), .B2(n21), .C(n20), .ZN(n31) );
  AOI221D0 U88 ( .A1(n25), .A2(search_data[20]), .B1(search_data[17]), .B2(n24), .C(n23), .ZN(n30) );
  AOI221D0 U89 ( .A1(n28), .A2(search_data[18]), .B1(search_data[15]), .B2(n27), .C(n26), .ZN(n29) );
  AOI221D0 U90 ( .A1(n35), .A2(search_data[0]), .B1(search_data[13]), .B2(n34), 
        .C(n33), .ZN(n48) );
  AOI221D0 U91 ( .A1(n38), .A2(search_data[14]), .B1(search_data[11]), .B2(n37), .C(n36), .ZN(n47) );
  AOI221D0 U92 ( .A1(n41), .A2(search_data[12]), .B1(search_data[9]), .B2(n40), 
        .C(n39), .ZN(n46) );
  AOI221D0 U93 ( .A1(n44), .A2(search_data[10]), .B1(search_data[25]), .B2(n43), .C(n42), .ZN(n45) );
  AOI221D0 U94 ( .A1(n51), .A2(search_data[7]), .B1(search_data[5]), .B2(n50), 
        .C(n49), .ZN(n65) );
  AOI221D0 U95 ( .A1(n54), .A2(search_data[16]), .B1(search_data[2]), .B2(n53), 
        .C(n52), .ZN(n64) );
  OAI221D0 U96 ( .A1(n57), .A2(search_data[3]), .B1(n56), .B2(search_data[6]), 
        .C(n55), .ZN(n62) );
  OAI221D0 U97 ( .A1(n60), .A2(search_data[1]), .B1(n59), .B2(search_data[4]), 
        .C(n58), .ZN(n61) );
  AO22D0 U98 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U99 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U100 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U101 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U102 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U103 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U104 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U105 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U106 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U107 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U108 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_28 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AN3D0 U4 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results) );
  ND4D0 U5 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  AO21D0 U6 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U7 ( .A1(reset), .A2(n70), .ZN(n71) );
  CKND2D1 U8 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  AOI21D2 U9 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  OAI22D0 U10 ( .A1(n19), .A2(search_data[8]), .B1(n18), .B2(search_data[21]), 
        .ZN(n17) );
  OAI22D0 U11 ( .A1(n12), .A2(search_data[26]), .B1(n11), .B2(search_data[23]), 
        .ZN(n10) );
  OAI22D0 U12 ( .A1(n9), .A2(search_data[28]), .B1(n8), .B2(search_data[24]), 
        .ZN(n7) );
  OAI22D0 U13 ( .A1(n6), .A2(search_data[30]), .B1(n5), .B2(search_data[27]), 
        .ZN(n4) );
  OAI22D0 U14 ( .A1(n3), .A2(search_data[31]), .B1(n2), .B2(search_data[29]), 
        .ZN(n1) );
  OAI22D0 U15 ( .A1(n22), .A2(search_data[22]), .B1(n21), .B2(search_data[19]), 
        .ZN(n20) );
  AOI22D0 U16 ( .A1(search_data[1]), .A2(n60), .B1(search_data[4]), .B2(n59), 
        .ZN(n58) );
  AOI22D0 U17 ( .A1(search_data[3]), .A2(n57), .B1(search_data[6]), .B2(n56), 
        .ZN(n55) );
  OAI22D0 U18 ( .A1(n54), .A2(search_data[16]), .B1(n53), .B2(search_data[2]), 
        .ZN(n52) );
  OAI22D0 U19 ( .A1(n51), .A2(search_data[7]), .B1(n50), .B2(search_data[5]), 
        .ZN(n49) );
  OAI22D0 U20 ( .A1(n44), .A2(search_data[10]), .B1(n43), .B2(search_data[25]), 
        .ZN(n42) );
  OAI22D0 U21 ( .A1(n41), .A2(search_data[12]), .B1(n40), .B2(search_data[9]), 
        .ZN(n39) );
  OAI22D0 U22 ( .A1(n38), .A2(search_data[14]), .B1(n37), .B2(search_data[11]), 
        .ZN(n36) );
  OAI22D0 U23 ( .A1(n35), .A2(search_data[0]), .B1(n34), .B2(search_data[13]), 
        .ZN(n33) );
  OAI22D0 U24 ( .A1(n28), .A2(search_data[18]), .B1(n27), .B2(search_data[15]), 
        .ZN(n26) );
  OAI22D0 U25 ( .A1(n25), .A2(search_data[20]), .B1(n24), .B2(search_data[17]), 
        .ZN(n23) );
  CKND0 U26 ( .I(read_value[10]), .ZN(n44) );
  CKND0 U27 ( .I(read_value[9]), .ZN(n40) );
  CKND0 U28 ( .I(read_value[12]), .ZN(n41) );
  CKND0 U29 ( .I(read_value[11]), .ZN(n37) );
  CKND0 U30 ( .I(read_value[14]), .ZN(n38) );
  CKND0 U31 ( .I(read_value[13]), .ZN(n34) );
  CKND0 U32 ( .I(read_value[0]), .ZN(n35) );
  CKND0 U33 ( .I(read_value[15]), .ZN(n27) );
  CKND0 U34 ( .I(read_value[18]), .ZN(n28) );
  CKND0 U35 ( .I(read_value[17]), .ZN(n24) );
  CKND0 U36 ( .I(read_value[20]), .ZN(n25) );
  CKND0 U37 ( .I(read_value[19]), .ZN(n21) );
  CKND0 U38 ( .I(read_value[22]), .ZN(n22) );
  CKND0 U39 ( .I(read_value[21]), .ZN(n18) );
  CKND0 U40 ( .I(read_value[8]), .ZN(n19) );
  CKND0 U41 ( .I(read_value[23]), .ZN(n11) );
  CKND0 U42 ( .I(read_value[26]), .ZN(n12) );
  CKND0 U43 ( .I(read_value[24]), .ZN(n8) );
  CKND0 U44 ( .I(read_value[28]), .ZN(n9) );
  CKND0 U45 ( .I(read_value[27]), .ZN(n5) );
  CKND0 U46 ( .I(read_value[30]), .ZN(n6) );
  CKND0 U47 ( .I(read_value[29]), .ZN(n2) );
  CKND0 U48 ( .I(read_value[31]), .ZN(n3) );
  CKND0 U49 ( .I(read_value[4]), .ZN(n59) );
  CKND0 U50 ( .I(read_value[1]), .ZN(n60) );
  CKND0 U51 ( .I(read_value[6]), .ZN(n56) );
  CKND0 U52 ( .I(read_value[3]), .ZN(n57) );
  CKND0 U53 ( .I(read_value[2]), .ZN(n53) );
  CKND0 U54 ( .I(read_value[16]), .ZN(n54) );
  CKND0 U55 ( .I(read_value[5]), .ZN(n50) );
  CKND0 U56 ( .I(read_value[7]), .ZN(n51) );
  CKND0 U57 ( .I(read_value[25]), .ZN(n43) );
  AO22D0 U58 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U59 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U60 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U61 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U62 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U63 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U64 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U65 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U66 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U67 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U68 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U69 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U70 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U71 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U72 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U73 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U74 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U75 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U76 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U77 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  NR2D1 U78 ( .A1(n62), .A2(n61), .ZN(n63) );
  ND4D1 U79 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .ZN(n67) );
  ND4D1 U80 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .ZN(n68) );
  ND4D1 U81 ( .A1(n16), .A2(n15), .A3(n14), .A4(n13), .ZN(n69) );
  AOI221D0 U82 ( .A1(n3), .A2(search_data[31]), .B1(search_data[29]), .B2(n2), 
        .C(n1), .ZN(n16) );
  AOI221D0 U83 ( .A1(n6), .A2(search_data[30]), .B1(search_data[27]), .B2(n5), 
        .C(n4), .ZN(n15) );
  AOI221D0 U84 ( .A1(n9), .A2(search_data[28]), .B1(search_data[24]), .B2(n8), 
        .C(n7), .ZN(n14) );
  AOI221D0 U85 ( .A1(n12), .A2(search_data[26]), .B1(search_data[23]), .B2(n11), .C(n10), .ZN(n13) );
  AOI221D0 U86 ( .A1(n19), .A2(search_data[8]), .B1(search_data[21]), .B2(n18), 
        .C(n17), .ZN(n32) );
  AOI221D0 U87 ( .A1(n22), .A2(search_data[22]), .B1(search_data[19]), .B2(n21), .C(n20), .ZN(n31) );
  AOI221D0 U88 ( .A1(n25), .A2(search_data[20]), .B1(search_data[17]), .B2(n24), .C(n23), .ZN(n30) );
  AOI221D0 U89 ( .A1(n28), .A2(search_data[18]), .B1(search_data[15]), .B2(n27), .C(n26), .ZN(n29) );
  AOI221D0 U90 ( .A1(n35), .A2(search_data[0]), .B1(search_data[13]), .B2(n34), 
        .C(n33), .ZN(n48) );
  AOI221D0 U91 ( .A1(n38), .A2(search_data[14]), .B1(search_data[11]), .B2(n37), .C(n36), .ZN(n47) );
  AOI221D0 U92 ( .A1(n41), .A2(search_data[12]), .B1(search_data[9]), .B2(n40), 
        .C(n39), .ZN(n46) );
  AOI221D0 U93 ( .A1(n44), .A2(search_data[10]), .B1(search_data[25]), .B2(n43), .C(n42), .ZN(n45) );
  AOI221D0 U94 ( .A1(n51), .A2(search_data[7]), .B1(search_data[5]), .B2(n50), 
        .C(n49), .ZN(n65) );
  AOI221D0 U95 ( .A1(n54), .A2(search_data[16]), .B1(search_data[2]), .B2(n53), 
        .C(n52), .ZN(n64) );
  OAI221D0 U96 ( .A1(n57), .A2(search_data[3]), .B1(n56), .B2(search_data[6]), 
        .C(n55), .ZN(n62) );
  OAI221D0 U97 ( .A1(n60), .A2(search_data[1]), .B1(n59), .B2(search_data[4]), 
        .C(n58), .ZN(n61) );
  AO22D0 U98 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U99 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U100 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), 
        .Z(data_i[2]) );
  AO22D0 U101 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), 
        .Z(data_i[3]) );
  AO22D0 U102 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), 
        .Z(data_i[4]) );
  AO22D0 U103 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), 
        .Z(data_i[5]) );
  AO22D0 U104 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), 
        .Z(data_i[6]) );
  AO22D0 U105 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U106 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U107 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U108 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_29 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AN3D0 U4 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results) );
  ND4D0 U5 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  AO21D0 U6 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U7 ( .A1(reset), .A2(n70), .ZN(n71) );
  CKND2D1 U8 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  AOI21D2 U9 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  AOI22D0 U10 ( .A1(search_data[1]), .A2(n60), .B1(search_data[4]), .B2(n59), 
        .ZN(n58) );
  AOI22D0 U11 ( .A1(search_data[3]), .A2(n57), .B1(search_data[6]), .B2(n56), 
        .ZN(n55) );
  OAI22D0 U12 ( .A1(n54), .A2(search_data[16]), .B1(n53), .B2(search_data[2]), 
        .ZN(n52) );
  OAI22D0 U13 ( .A1(n51), .A2(search_data[7]), .B1(n50), .B2(search_data[5]), 
        .ZN(n49) );
  OAI22D0 U14 ( .A1(n44), .A2(search_data[10]), .B1(n43), .B2(search_data[25]), 
        .ZN(n42) );
  OAI22D0 U15 ( .A1(n41), .A2(search_data[12]), .B1(n40), .B2(search_data[9]), 
        .ZN(n39) );
  OAI22D0 U16 ( .A1(n38), .A2(search_data[14]), .B1(n37), .B2(search_data[11]), 
        .ZN(n36) );
  OAI22D0 U17 ( .A1(n35), .A2(search_data[0]), .B1(n34), .B2(search_data[13]), 
        .ZN(n33) );
  OAI22D0 U18 ( .A1(n28), .A2(search_data[18]), .B1(n27), .B2(search_data[15]), 
        .ZN(n26) );
  OAI22D0 U19 ( .A1(n25), .A2(search_data[20]), .B1(n24), .B2(search_data[17]), 
        .ZN(n23) );
  OAI22D0 U20 ( .A1(n22), .A2(search_data[22]), .B1(n21), .B2(search_data[19]), 
        .ZN(n20) );
  OAI22D0 U21 ( .A1(n19), .A2(search_data[8]), .B1(n18), .B2(search_data[21]), 
        .ZN(n17) );
  OAI22D0 U22 ( .A1(n12), .A2(search_data[26]), .B1(n11), .B2(search_data[23]), 
        .ZN(n10) );
  OAI22D0 U23 ( .A1(n9), .A2(search_data[28]), .B1(n8), .B2(search_data[24]), 
        .ZN(n7) );
  OAI22D0 U24 ( .A1(n6), .A2(search_data[30]), .B1(n5), .B2(search_data[27]), 
        .ZN(n4) );
  OAI22D0 U25 ( .A1(n3), .A2(search_data[31]), .B1(n2), .B2(search_data[29]), 
        .ZN(n1) );
  CKND0 U26 ( .I(read_value[15]), .ZN(n27) );
  CKND0 U27 ( .I(read_value[18]), .ZN(n28) );
  CKND0 U28 ( .I(read_value[17]), .ZN(n24) );
  CKND0 U29 ( .I(read_value[20]), .ZN(n25) );
  CKND0 U30 ( .I(read_value[19]), .ZN(n21) );
  CKND0 U31 ( .I(read_value[22]), .ZN(n22) );
  CKND0 U32 ( .I(read_value[21]), .ZN(n18) );
  CKND0 U33 ( .I(read_value[8]), .ZN(n19) );
  CKND0 U34 ( .I(read_value[23]), .ZN(n11) );
  CKND0 U35 ( .I(read_value[26]), .ZN(n12) );
  CKND0 U36 ( .I(read_value[24]), .ZN(n8) );
  CKND0 U37 ( .I(read_value[28]), .ZN(n9) );
  CKND0 U38 ( .I(read_value[27]), .ZN(n5) );
  CKND0 U39 ( .I(read_value[30]), .ZN(n6) );
  CKND0 U40 ( .I(read_value[29]), .ZN(n2) );
  CKND0 U41 ( .I(read_value[31]), .ZN(n3) );
  CKND0 U42 ( .I(read_value[4]), .ZN(n59) );
  CKND0 U43 ( .I(read_value[10]), .ZN(n44) );
  CKND0 U44 ( .I(read_value[25]), .ZN(n43) );
  CKND0 U45 ( .I(read_value[9]), .ZN(n40) );
  CKND0 U46 ( .I(read_value[12]), .ZN(n41) );
  CKND0 U47 ( .I(read_value[7]), .ZN(n51) );
  CKND0 U48 ( .I(read_value[5]), .ZN(n50) );
  CKND0 U49 ( .I(read_value[11]), .ZN(n37) );
  CKND0 U50 ( .I(read_value[16]), .ZN(n54) );
  CKND0 U51 ( .I(read_value[2]), .ZN(n53) );
  CKND0 U52 ( .I(read_value[0]), .ZN(n35) );
  CKND0 U53 ( .I(read_value[1]), .ZN(n60) );
  CKND0 U54 ( .I(read_value[14]), .ZN(n38) );
  CKND0 U55 ( .I(read_value[6]), .ZN(n56) );
  CKND0 U56 ( .I(read_value[3]), .ZN(n57) );
  CKND0 U57 ( .I(read_value[13]), .ZN(n34) );
  AO22D0 U58 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U59 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U60 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U61 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U62 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U63 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U64 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U65 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U66 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U67 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U68 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U69 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U70 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U71 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U72 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U73 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U74 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  AO22D0 U75 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U76 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U77 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  NR2D1 U78 ( .A1(n62), .A2(n61), .ZN(n63) );
  ND4D1 U79 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .ZN(n67) );
  ND4D1 U80 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .ZN(n68) );
  ND4D1 U81 ( .A1(n16), .A2(n15), .A3(n14), .A4(n13), .ZN(n69) );
  AOI221D0 U82 ( .A1(n3), .A2(search_data[31]), .B1(search_data[29]), .B2(n2), 
        .C(n1), .ZN(n16) );
  AOI221D0 U83 ( .A1(n6), .A2(search_data[30]), .B1(search_data[27]), .B2(n5), 
        .C(n4), .ZN(n15) );
  AOI221D0 U84 ( .A1(n9), .A2(search_data[28]), .B1(search_data[24]), .B2(n8), 
        .C(n7), .ZN(n14) );
  AOI221D0 U85 ( .A1(n12), .A2(search_data[26]), .B1(search_data[23]), .B2(n11), .C(n10), .ZN(n13) );
  AOI221D0 U86 ( .A1(n19), .A2(search_data[8]), .B1(search_data[21]), .B2(n18), 
        .C(n17), .ZN(n32) );
  AOI221D0 U87 ( .A1(n22), .A2(search_data[22]), .B1(search_data[19]), .B2(n21), .C(n20), .ZN(n31) );
  AOI221D0 U88 ( .A1(n25), .A2(search_data[20]), .B1(search_data[17]), .B2(n24), .C(n23), .ZN(n30) );
  AOI221D0 U89 ( .A1(n28), .A2(search_data[18]), .B1(search_data[15]), .B2(n27), .C(n26), .ZN(n29) );
  AOI221D0 U90 ( .A1(n35), .A2(search_data[0]), .B1(search_data[13]), .B2(n34), 
        .C(n33), .ZN(n48) );
  AOI221D0 U91 ( .A1(n38), .A2(search_data[14]), .B1(search_data[11]), .B2(n37), .C(n36), .ZN(n47) );
  AOI221D0 U92 ( .A1(n41), .A2(search_data[12]), .B1(search_data[9]), .B2(n40), 
        .C(n39), .ZN(n46) );
  AOI221D0 U93 ( .A1(n44), .A2(search_data[10]), .B1(search_data[25]), .B2(n43), .C(n42), .ZN(n45) );
  AOI221D0 U94 ( .A1(n51), .A2(search_data[7]), .B1(search_data[5]), .B2(n50), 
        .C(n49), .ZN(n65) );
  AOI221D0 U95 ( .A1(n54), .A2(search_data[16]), .B1(search_data[2]), .B2(n53), 
        .C(n52), .ZN(n64) );
  OAI221D0 U96 ( .A1(n57), .A2(search_data[3]), .B1(n56), .B2(search_data[6]), 
        .C(n55), .ZN(n62) );
  OAI221D0 U97 ( .A1(n60), .A2(search_data[1]), .B1(n59), .B2(search_data[4]), 
        .C(n58), .ZN(n61) );
  AO22D0 U98 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U99 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U100 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), 
        .Z(data_i[2]) );
  AO22D0 U101 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), 
        .Z(data_i[3]) );
  AO22D0 U102 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), 
        .Z(data_i[4]) );
  AO22D0 U103 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), 
        .Z(data_i[5]) );
  AO22D0 U104 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), 
        .Z(data_i[6]) );
  AO22D0 U105 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U106 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U107 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U108 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_30 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AN3D0 U4 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results) );
  AO21D0 U5 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  ND4D0 U6 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  NR2D2 U7 ( .A1(reset), .A2(n70), .ZN(n71) );
  CKND2D1 U8 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  AOI21D2 U9 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  AOI22D0 U10 ( .A1(search_data[1]), .A2(n60), .B1(search_data[4]), .B2(n59), 
        .ZN(n58) );
  AOI22D0 U11 ( .A1(search_data[3]), .A2(n57), .B1(search_data[6]), .B2(n56), 
        .ZN(n55) );
  OAI22D0 U12 ( .A1(n54), .A2(search_data[16]), .B1(n53), .B2(search_data[2]), 
        .ZN(n52) );
  OAI22D0 U13 ( .A1(n51), .A2(search_data[7]), .B1(n50), .B2(search_data[5]), 
        .ZN(n49) );
  OAI22D0 U14 ( .A1(n44), .A2(search_data[10]), .B1(n43), .B2(search_data[25]), 
        .ZN(n42) );
  OAI22D0 U15 ( .A1(n41), .A2(search_data[12]), .B1(n40), .B2(search_data[9]), 
        .ZN(n39) );
  OAI22D0 U16 ( .A1(n38), .A2(search_data[14]), .B1(n37), .B2(search_data[11]), 
        .ZN(n36) );
  OAI22D0 U17 ( .A1(n35), .A2(search_data[0]), .B1(n34), .B2(search_data[13]), 
        .ZN(n33) );
  OAI22D0 U18 ( .A1(n28), .A2(search_data[18]), .B1(n27), .B2(search_data[15]), 
        .ZN(n26) );
  OAI22D0 U19 ( .A1(n25), .A2(search_data[20]), .B1(n24), .B2(search_data[17]), 
        .ZN(n23) );
  OAI22D0 U20 ( .A1(n22), .A2(search_data[22]), .B1(n21), .B2(search_data[19]), 
        .ZN(n20) );
  OAI22D0 U21 ( .A1(n19), .A2(search_data[8]), .B1(n18), .B2(search_data[21]), 
        .ZN(n17) );
  OAI22D0 U22 ( .A1(n12), .A2(search_data[26]), .B1(n11), .B2(search_data[23]), 
        .ZN(n10) );
  OAI22D0 U23 ( .A1(n9), .A2(search_data[28]), .B1(n8), .B2(search_data[24]), 
        .ZN(n7) );
  OAI22D0 U24 ( .A1(n6), .A2(search_data[30]), .B1(n5), .B2(search_data[27]), 
        .ZN(n4) );
  OAI22D0 U25 ( .A1(n3), .A2(search_data[31]), .B1(n2), .B2(search_data[29]), 
        .ZN(n1) );
  CKND0 U26 ( .I(read_value[31]), .ZN(n3) );
  CKND0 U27 ( .I(read_value[29]), .ZN(n2) );
  CKND0 U28 ( .I(read_value[30]), .ZN(n6) );
  CKND0 U29 ( .I(read_value[27]), .ZN(n5) );
  CKND0 U30 ( .I(read_value[28]), .ZN(n9) );
  CKND0 U31 ( .I(read_value[24]), .ZN(n8) );
  CKND0 U32 ( .I(read_value[26]), .ZN(n12) );
  CKND0 U33 ( .I(read_value[23]), .ZN(n11) );
  CKND0 U34 ( .I(read_value[8]), .ZN(n19) );
  CKND0 U35 ( .I(read_value[21]), .ZN(n18) );
  CKND0 U36 ( .I(read_value[22]), .ZN(n22) );
  CKND0 U37 ( .I(read_value[19]), .ZN(n21) );
  CKND0 U38 ( .I(read_value[4]), .ZN(n59) );
  CKND0 U39 ( .I(read_value[20]), .ZN(n25) );
  CKND0 U40 ( .I(read_value[17]), .ZN(n24) );
  CKND0 U41 ( .I(read_value[1]), .ZN(n60) );
  CKND0 U42 ( .I(read_value[18]), .ZN(n28) );
  CKND0 U43 ( .I(read_value[15]), .ZN(n27) );
  CKND0 U44 ( .I(read_value[6]), .ZN(n56) );
  CKND0 U45 ( .I(read_value[3]), .ZN(n57) );
  CKND0 U46 ( .I(read_value[0]), .ZN(n35) );
  CKND0 U47 ( .I(read_value[13]), .ZN(n34) );
  CKND0 U48 ( .I(read_value[2]), .ZN(n53) );
  CKND0 U49 ( .I(read_value[14]), .ZN(n38) );
  CKND0 U50 ( .I(read_value[16]), .ZN(n54) );
  CKND0 U51 ( .I(read_value[11]), .ZN(n37) );
  CKND0 U52 ( .I(read_value[12]), .ZN(n41) );
  CKND0 U53 ( .I(read_value[9]), .ZN(n40) );
  CKND0 U54 ( .I(read_value[5]), .ZN(n50) );
  CKND0 U55 ( .I(read_value[10]), .ZN(n44) );
  CKND0 U56 ( .I(read_value[25]), .ZN(n43) );
  CKND0 U57 ( .I(read_value[7]), .ZN(n51) );
  AO22D0 U58 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U59 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U60 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U61 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U62 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U63 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U64 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U65 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U66 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U67 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U68 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U69 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U70 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U71 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U72 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U73 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U74 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U75 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U76 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U77 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  NR2D1 U78 ( .A1(n62), .A2(n61), .ZN(n63) );
  ND4D1 U79 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .ZN(n67) );
  ND4D1 U80 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .ZN(n68) );
  ND4D1 U81 ( .A1(n16), .A2(n15), .A3(n14), .A4(n13), .ZN(n69) );
  AOI221D0 U82 ( .A1(n3), .A2(search_data[31]), .B1(search_data[29]), .B2(n2), 
        .C(n1), .ZN(n16) );
  AOI221D0 U83 ( .A1(n6), .A2(search_data[30]), .B1(search_data[27]), .B2(n5), 
        .C(n4), .ZN(n15) );
  AOI221D0 U84 ( .A1(n9), .A2(search_data[28]), .B1(search_data[24]), .B2(n8), 
        .C(n7), .ZN(n14) );
  AOI221D0 U85 ( .A1(n12), .A2(search_data[26]), .B1(search_data[23]), .B2(n11), .C(n10), .ZN(n13) );
  AOI221D0 U86 ( .A1(n19), .A2(search_data[8]), .B1(search_data[21]), .B2(n18), 
        .C(n17), .ZN(n32) );
  AOI221D0 U87 ( .A1(n22), .A2(search_data[22]), .B1(search_data[19]), .B2(n21), .C(n20), .ZN(n31) );
  AOI221D0 U88 ( .A1(n25), .A2(search_data[20]), .B1(search_data[17]), .B2(n24), .C(n23), .ZN(n30) );
  AOI221D0 U89 ( .A1(n28), .A2(search_data[18]), .B1(search_data[15]), .B2(n27), .C(n26), .ZN(n29) );
  AOI221D0 U90 ( .A1(n35), .A2(search_data[0]), .B1(search_data[13]), .B2(n34), 
        .C(n33), .ZN(n48) );
  AOI221D0 U91 ( .A1(n38), .A2(search_data[14]), .B1(search_data[11]), .B2(n37), .C(n36), .ZN(n47) );
  AOI221D0 U92 ( .A1(n41), .A2(search_data[12]), .B1(search_data[9]), .B2(n40), 
        .C(n39), .ZN(n46) );
  AOI221D0 U93 ( .A1(n44), .A2(search_data[10]), .B1(search_data[25]), .B2(n43), .C(n42), .ZN(n45) );
  AOI221D0 U94 ( .A1(n51), .A2(search_data[7]), .B1(search_data[5]), .B2(n50), 
        .C(n49), .ZN(n65) );
  AOI221D0 U95 ( .A1(n54), .A2(search_data[16]), .B1(search_data[2]), .B2(n53), 
        .C(n52), .ZN(n64) );
  OAI221D0 U96 ( .A1(n57), .A2(search_data[3]), .B1(n56), .B2(search_data[6]), 
        .C(n55), .ZN(n62) );
  OAI221D0 U97 ( .A1(n60), .A2(search_data[1]), .B1(n59), .B2(search_data[4]), 
        .C(n58), .ZN(n61) );
  AO22D0 U98 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U99 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U100 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), 
        .Z(data_i[2]) );
  AO22D0 U101 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), 
        .Z(data_i[3]) );
  AO22D0 U102 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), 
        .Z(data_i[4]) );
  AO22D0 U103 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), 
        .Z(data_i[5]) );
  AO22D0 U104 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), 
        .Z(data_i[6]) );
  AO22D0 U105 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U106 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U107 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U108 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module cam_word_31 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   valid_i, valid_o, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72;
  wire   [31:0] data_i;

  DFQD1 \data_ff/data_reg[0]  ( .D(data_i[0]), .CP(clk), .Q(read_value[0]) );
  DFQD1 \data_ff/data_reg[1]  ( .D(data_i[1]), .CP(clk), .Q(read_value[1]) );
  DFQD1 \data_ff/data_reg[2]  ( .D(data_i[2]), .CP(clk), .Q(read_value[2]) );
  DFQD1 \data_ff/data_reg[3]  ( .D(data_i[3]), .CP(clk), .Q(read_value[3]) );
  DFQD1 \data_ff/data_reg[4]  ( .D(data_i[4]), .CP(clk), .Q(read_value[4]) );
  DFQD1 \data_ff/data_reg[5]  ( .D(data_i[5]), .CP(clk), .Q(read_value[5]) );
  DFQD1 \data_ff/data_reg[6]  ( .D(data_i[6]), .CP(clk), .Q(read_value[6]) );
  DFQD1 \data_ff/data_reg[7]  ( .D(data_i[7]), .CP(clk), .Q(read_value[7]) );
  DFQD1 \data_ff/data_reg[8]  ( .D(data_i[8]), .CP(clk), .Q(read_value[8]) );
  DFQD1 \data_ff/data_reg[9]  ( .D(data_i[9]), .CP(clk), .Q(read_value[9]) );
  DFQD1 \data_ff/data_reg[10]  ( .D(data_i[10]), .CP(clk), .Q(read_value[10])
         );
  DFQD1 \data_ff/data_reg[11]  ( .D(data_i[11]), .CP(clk), .Q(read_value[11])
         );
  DFQD1 \data_ff/data_reg[12]  ( .D(data_i[12]), .CP(clk), .Q(read_value[12])
         );
  DFQD1 \data_ff/data_reg[13]  ( .D(data_i[13]), .CP(clk), .Q(read_value[13])
         );
  DFQD1 \data_ff/data_reg[14]  ( .D(data_i[14]), .CP(clk), .Q(read_value[14])
         );
  DFQD1 \data_ff/data_reg[15]  ( .D(data_i[15]), .CP(clk), .Q(read_value[15])
         );
  DFQD1 \data_ff/data_reg[16]  ( .D(data_i[16]), .CP(clk), .Q(read_value[16])
         );
  DFQD1 \data_ff/data_reg[17]  ( .D(data_i[17]), .CP(clk), .Q(read_value[17])
         );
  DFQD1 \data_ff/data_reg[18]  ( .D(data_i[18]), .CP(clk), .Q(read_value[18])
         );
  DFQD1 \data_ff/data_reg[19]  ( .D(data_i[19]), .CP(clk), .Q(read_value[19])
         );
  DFQD1 \data_ff/data_reg[20]  ( .D(data_i[20]), .CP(clk), .Q(read_value[20])
         );
  DFQD1 \data_ff/data_reg[21]  ( .D(data_i[21]), .CP(clk), .Q(read_value[21])
         );
  DFQD1 \data_ff/data_reg[22]  ( .D(data_i[22]), .CP(clk), .Q(read_value[22])
         );
  DFQD1 \data_ff/data_reg[23]  ( .D(data_i[23]), .CP(clk), .Q(read_value[23])
         );
  DFQD1 \data_ff/data_reg[24]  ( .D(data_i[24]), .CP(clk), .Q(read_value[24])
         );
  DFQD1 \data_ff/data_reg[25]  ( .D(data_i[25]), .CP(clk), .Q(read_value[25])
         );
  DFQD1 \data_ff/data_reg[26]  ( .D(data_i[26]), .CP(clk), .Q(read_value[26])
         );
  DFQD1 \data_ff/data_reg[27]  ( .D(data_i[27]), .CP(clk), .Q(read_value[27])
         );
  DFQD1 \data_ff/data_reg[28]  ( .D(data_i[28]), .CP(clk), .Q(read_value[28])
         );
  DFQD1 \data_ff/data_reg[29]  ( .D(data_i[29]), .CP(clk), .Q(read_value[29])
         );
  DFQD1 \data_ff/data_reg[30]  ( .D(data_i[30]), .CP(clk), .Q(read_value[30])
         );
  DFQD1 \data_ff/data_reg[31]  ( .D(data_i[31]), .CP(clk), .Q(read_value[31])
         );
  DFQD1 \valid_ff/data_reg[0]  ( .D(valid_i), .CP(clk), .Q(valid_o) );
  NR4D0 U3 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(search_results) );
  AN3D0 U4 ( .A1(valid_o), .A2(dec_read_index), .A3(read), .Z(read_results) );
  ND4D0 U5 ( .A1(n65), .A2(search), .A3(n64), .A4(n63), .ZN(n66) );
  AO21D0 U6 ( .A1(n72), .A2(valid_o), .B(n71), .Z(valid_i) );
  NR2D2 U7 ( .A1(reset), .A2(n70), .ZN(n71) );
  OAI22D0 U8 ( .A1(n25), .A2(search_data[20]), .B1(n24), .B2(search_data[17]), 
        .ZN(n23) );
  OAI22D0 U9 ( .A1(n22), .A2(search_data[22]), .B1(n21), .B2(search_data[19]), 
        .ZN(n20) );
  OAI22D0 U10 ( .A1(n19), .A2(search_data[8]), .B1(n18), .B2(search_data[21]), 
        .ZN(n17) );
  OAI22D0 U11 ( .A1(n41), .A2(search_data[12]), .B1(n40), .B2(search_data[9]), 
        .ZN(n39) );
  OAI22D0 U12 ( .A1(n35), .A2(search_data[0]), .B1(n34), .B2(search_data[13]), 
        .ZN(n33) );
  OAI22D0 U13 ( .A1(n38), .A2(search_data[14]), .B1(n37), .B2(search_data[11]), 
        .ZN(n36) );
  OAI22D0 U14 ( .A1(n28), .A2(search_data[18]), .B1(n27), .B2(search_data[15]), 
        .ZN(n26) );
  OAI22D0 U15 ( .A1(n12), .A2(search_data[26]), .B1(n11), .B2(search_data[23]), 
        .ZN(n10) );
  OAI22D0 U16 ( .A1(n9), .A2(search_data[28]), .B1(n8), .B2(search_data[24]), 
        .ZN(n7) );
  OAI22D0 U17 ( .A1(n6), .A2(search_data[30]), .B1(n5), .B2(search_data[27]), 
        .ZN(n4) );
  OAI22D0 U18 ( .A1(n3), .A2(search_data[31]), .B1(n2), .B2(search_data[29]), 
        .ZN(n1) );
  AOI22D0 U19 ( .A1(search_data[1]), .A2(n60), .B1(search_data[4]), .B2(n59), 
        .ZN(n58) );
  AOI22D0 U20 ( .A1(search_data[3]), .A2(n57), .B1(search_data[6]), .B2(n56), 
        .ZN(n55) );
  OAI22D0 U21 ( .A1(n54), .A2(search_data[16]), .B1(n53), .B2(search_data[2]), 
        .ZN(n52) );
  OAI22D0 U22 ( .A1(n51), .A2(search_data[7]), .B1(n50), .B2(search_data[5]), 
        .ZN(n49) );
  OAI22D0 U23 ( .A1(n44), .A2(search_data[10]), .B1(n43), .B2(search_data[25]), 
        .ZN(n42) );
  AOI21D2 U24 ( .A1(write), .A2(dec_write_index), .B(reset), .ZN(n72) );
  CKND2D1 U25 ( .A1(write), .A2(dec_write_index), .ZN(n70) );
  CKND0 U26 ( .I(read_value[12]), .ZN(n41) );
  CKND0 U27 ( .I(read_value[11]), .ZN(n37) );
  CKND0 U28 ( .I(read_value[14]), .ZN(n38) );
  CKND0 U29 ( .I(read_value[7]), .ZN(n51) );
  CKND0 U30 ( .I(read_value[5]), .ZN(n50) );
  CKND0 U31 ( .I(read_value[16]), .ZN(n54) );
  CKND0 U32 ( .I(read_value[2]), .ZN(n53) );
  CKND0 U33 ( .I(read_value[3]), .ZN(n57) );
  CKND0 U34 ( .I(read_value[25]), .ZN(n43) );
  CKND0 U35 ( .I(read_value[6]), .ZN(n56) );
  CKND0 U36 ( .I(read_value[1]), .ZN(n60) );
  CKND0 U37 ( .I(read_value[4]), .ZN(n59) );
  CKND0 U38 ( .I(read_value[10]), .ZN(n44) );
  CKND0 U39 ( .I(read_value[9]), .ZN(n40) );
  CKND0 U40 ( .I(read_value[23]), .ZN(n11) );
  CKND0 U41 ( .I(read_value[26]), .ZN(n12) );
  CKND0 U42 ( .I(read_value[24]), .ZN(n8) );
  CKND0 U43 ( .I(read_value[28]), .ZN(n9) );
  CKND0 U44 ( .I(read_value[27]), .ZN(n5) );
  CKND0 U45 ( .I(read_value[30]), .ZN(n6) );
  CKND0 U46 ( .I(read_value[29]), .ZN(n2) );
  CKND0 U47 ( .I(read_value[31]), .ZN(n3) );
  CKND0 U48 ( .I(read_value[17]), .ZN(n24) );
  CKND0 U49 ( .I(read_value[20]), .ZN(n25) );
  CKND0 U50 ( .I(read_value[18]), .ZN(n28) );
  CKND0 U51 ( .I(read_value[19]), .ZN(n21) );
  CKND0 U52 ( .I(read_value[15]), .ZN(n27) );
  CKND0 U53 ( .I(read_value[22]), .ZN(n22) );
  CKND0 U54 ( .I(read_value[0]), .ZN(n35) );
  CKND0 U55 ( .I(read_value[21]), .ZN(n18) );
  CKND0 U56 ( .I(read_value[8]), .ZN(n19) );
  CKND0 U57 ( .I(read_value[13]), .ZN(n34) );
  AO22D0 U58 ( .A1(read_value[25]), .A2(n72), .B1(n71), .B2(write_data[25]), 
        .Z(data_i[25]) );
  AO22D0 U59 ( .A1(read_value[13]), .A2(n72), .B1(n71), .B2(write_data[13]), 
        .Z(data_i[13]) );
  AO22D0 U60 ( .A1(read_value[12]), .A2(n72), .B1(n71), .B2(write_data[12]), 
        .Z(data_i[12]) );
  AO22D0 U61 ( .A1(read_value[11]), .A2(n72), .B1(n71), .B2(write_data[11]), 
        .Z(data_i[11]) );
  AO22D0 U62 ( .A1(read_value[10]), .A2(n72), .B1(n71), .B2(write_data[10]), 
        .Z(data_i[10]) );
  AO22D0 U63 ( .A1(read_value[9]), .A2(n72), .B1(n71), .B2(write_data[9]), .Z(
        data_i[9]) );
  AO22D0 U64 ( .A1(read_value[8]), .A2(n72), .B1(n71), .B2(write_data[8]), .Z(
        data_i[8]) );
  AO22D0 U65 ( .A1(read_value[7]), .A2(n72), .B1(n71), .B2(write_data[7]), .Z(
        data_i[7]) );
  AO22D0 U66 ( .A1(read_value[24]), .A2(n72), .B1(n71), .B2(write_data[24]), 
        .Z(data_i[24]) );
  AO22D0 U67 ( .A1(read_value[23]), .A2(n72), .B1(n71), .B2(write_data[23]), 
        .Z(data_i[23]) );
  AO22D0 U68 ( .A1(read_value[22]), .A2(n72), .B1(n71), .B2(write_data[22]), 
        .Z(data_i[22]) );
  AO22D0 U69 ( .A1(read_value[21]), .A2(n72), .B1(n71), .B2(write_data[21]), 
        .Z(data_i[21]) );
  AO22D0 U70 ( .A1(read_value[20]), .A2(n72), .B1(n71), .B2(write_data[20]), 
        .Z(data_i[20]) );
  AO22D0 U71 ( .A1(read_value[19]), .A2(n72), .B1(n71), .B2(write_data[19]), 
        .Z(data_i[19]) );
  AO22D0 U72 ( .A1(read_value[18]), .A2(n72), .B1(n71), .B2(write_data[18]), 
        .Z(data_i[18]) );
  AO22D0 U73 ( .A1(read_value[17]), .A2(n72), .B1(n71), .B2(write_data[17]), 
        .Z(data_i[17]) );
  AO22D0 U74 ( .A1(read_value[16]), .A2(n72), .B1(n71), .B2(write_data[16]), 
        .Z(data_i[16]) );
  AO22D0 U75 ( .A1(read_value[15]), .A2(n72), .B1(n71), .B2(write_data[15]), 
        .Z(data_i[15]) );
  AO22D0 U76 ( .A1(read_value[14]), .A2(n72), .B1(n71), .B2(write_data[14]), 
        .Z(data_i[14]) );
  AO22D0 U77 ( .A1(read_value[26]), .A2(n72), .B1(n71), .B2(write_data[26]), 
        .Z(data_i[26]) );
  NR2D1 U78 ( .A1(n62), .A2(n61), .ZN(n63) );
  ND4D1 U79 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .ZN(n67) );
  ND4D1 U80 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .ZN(n68) );
  ND4D1 U81 ( .A1(n16), .A2(n15), .A3(n14), .A4(n13), .ZN(n69) );
  AOI221D0 U82 ( .A1(n3), .A2(search_data[31]), .B1(search_data[29]), .B2(n2), 
        .C(n1), .ZN(n16) );
  AOI221D0 U83 ( .A1(n6), .A2(search_data[30]), .B1(search_data[27]), .B2(n5), 
        .C(n4), .ZN(n15) );
  AOI221D0 U84 ( .A1(n9), .A2(search_data[28]), .B1(search_data[24]), .B2(n8), 
        .C(n7), .ZN(n14) );
  AOI221D0 U85 ( .A1(n12), .A2(search_data[26]), .B1(search_data[23]), .B2(n11), .C(n10), .ZN(n13) );
  AOI221D0 U86 ( .A1(n19), .A2(search_data[8]), .B1(search_data[21]), .B2(n18), 
        .C(n17), .ZN(n32) );
  AOI221D0 U87 ( .A1(n22), .A2(search_data[22]), .B1(search_data[19]), .B2(n21), .C(n20), .ZN(n31) );
  AOI221D0 U88 ( .A1(n25), .A2(search_data[20]), .B1(search_data[17]), .B2(n24), .C(n23), .ZN(n30) );
  AOI221D0 U89 ( .A1(n28), .A2(search_data[18]), .B1(search_data[15]), .B2(n27), .C(n26), .ZN(n29) );
  AOI221D0 U90 ( .A1(n35), .A2(search_data[0]), .B1(search_data[13]), .B2(n34), 
        .C(n33), .ZN(n48) );
  AOI221D0 U91 ( .A1(n38), .A2(search_data[14]), .B1(search_data[11]), .B2(n37), .C(n36), .ZN(n47) );
  AOI221D0 U92 ( .A1(n41), .A2(search_data[12]), .B1(search_data[9]), .B2(n40), 
        .C(n39), .ZN(n46) );
  AOI221D0 U93 ( .A1(n44), .A2(search_data[10]), .B1(search_data[25]), .B2(n43), .C(n42), .ZN(n45) );
  AOI221D0 U94 ( .A1(n51), .A2(search_data[7]), .B1(search_data[5]), .B2(n50), 
        .C(n49), .ZN(n65) );
  AOI221D0 U95 ( .A1(n54), .A2(search_data[16]), .B1(search_data[2]), .B2(n53), 
        .C(n52), .ZN(n64) );
  OAI221D0 U96 ( .A1(n57), .A2(search_data[3]), .B1(n56), .B2(search_data[6]), 
        .C(n55), .ZN(n62) );
  OAI221D0 U97 ( .A1(n60), .A2(search_data[1]), .B1(n59), .B2(search_data[4]), 
        .C(n58), .ZN(n61) );
  AO22D0 U98 ( .A1(read_value[0]), .A2(n72), .B1(n71), .B2(write_data[0]), .Z(
        data_i[0]) );
  AO22D0 U99 ( .A1(read_value[1]), .A2(n72), .B1(n71), .B2(write_data[1]), .Z(
        data_i[1]) );
  AO22D0 U100 ( .A1(read_value[2]), .A2(n72), .B1(n71), .B2(write_data[2]), 
        .Z(data_i[2]) );
  AO22D0 U101 ( .A1(read_value[3]), .A2(n72), .B1(n71), .B2(write_data[3]), 
        .Z(data_i[3]) );
  AO22D0 U102 ( .A1(read_value[4]), .A2(n72), .B1(n71), .B2(write_data[4]), 
        .Z(data_i[4]) );
  AO22D0 U103 ( .A1(read_value[5]), .A2(n72), .B1(n71), .B2(write_data[5]), 
        .Z(data_i[5]) );
  AO22D0 U104 ( .A1(read_value[6]), .A2(n72), .B1(n71), .B2(write_data[6]), 
        .Z(data_i[6]) );
  AO22D0 U105 ( .A1(read_value[27]), .A2(n72), .B1(n71), .B2(write_data[27]), 
        .Z(data_i[27]) );
  AO22D0 U106 ( .A1(read_value[28]), .A2(n72), .B1(n71), .B2(write_data[28]), 
        .Z(data_i[28]) );
  AO22D0 U107 ( .A1(read_value[29]), .A2(n72), .B1(n71), .B2(write_data[29]), 
        .Z(data_i[29]) );
  AO22D0 U108 ( .A1(read_value[30]), .A2(n72), .B1(n71), .B2(write_data[30]), 
        .Z(data_i[30]) );
  AO22D0 U109 ( .A1(read_value[31]), .A2(n72), .B1(n71), .B2(write_data[31]), 
        .Z(data_i[31]) );
endmodule


module decoder_5_32_1 ( decoder_i, decoder_o );
  input [4:0] decoder_i;
  output [31:0] decoder_o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;

  ND2D1 U1 ( .A1(n2), .A2(n1), .ZN(n18) );
  NR2D0 U2 ( .A1(n11), .A2(n17), .ZN(decoder_o[12]) );
  NR2D0 U3 ( .A1(n11), .A2(n15), .ZN(decoder_o[14]) );
  NR2D0 U4 ( .A1(n12), .A2(n17), .ZN(decoder_o[8]) );
  NR2D0 U5 ( .A1(n12), .A2(n16), .ZN(decoder_o[9]) );
  NR2D0 U6 ( .A1(n12), .A2(n15), .ZN(decoder_o[10]) );
  NR2D0 U7 ( .A1(n12), .A2(n14), .ZN(decoder_o[11]) );
  NR2D0 U8 ( .A1(n13), .A2(n17), .ZN(decoder_o[4]) );
  NR2D0 U9 ( .A1(n13), .A2(n16), .ZN(decoder_o[5]) );
  NR2D0 U10 ( .A1(n13), .A2(n15), .ZN(decoder_o[6]) );
  NR2D0 U11 ( .A1(n13), .A2(n14), .ZN(decoder_o[7]) );
  NR2D0 U12 ( .A1(n18), .A2(n17), .ZN(decoder_o[0]) );
  NR2D0 U13 ( .A1(n18), .A2(n16), .ZN(decoder_o[1]) );
  NR2D0 U14 ( .A1(n18), .A2(n15), .ZN(decoder_o[2]) );
  NR2D0 U15 ( .A1(n18), .A2(n14), .ZN(decoder_o[3]) );
  NR2XD0 U16 ( .A1(n4), .A2(n18), .ZN(decoder_o[18]) );
  NR2D0 U17 ( .A1(n4), .A2(n13), .ZN(decoder_o[22]) );
  NR2D0 U18 ( .A1(n4), .A2(n12), .ZN(decoder_o[26]) );
  NR2D0 U19 ( .A1(n11), .A2(n4), .ZN(decoder_o[30]) );
  NR2D0 U20 ( .A1(n11), .A2(n6), .ZN(decoder_o[28]) );
  NR2D0 U21 ( .A1(n3), .A2(n13), .ZN(decoder_o[23]) );
  NR2D0 U22 ( .A1(n5), .A2(n13), .ZN(decoder_o[21]) );
  NR2D0 U23 ( .A1(n6), .A2(n13), .ZN(decoder_o[20]) );
  NR2D0 U24 ( .A1(n3), .A2(n12), .ZN(decoder_o[27]) );
  NR2D0 U25 ( .A1(n5), .A2(n12), .ZN(decoder_o[25]) );
  NR2D0 U26 ( .A1(n6), .A2(n12), .ZN(decoder_o[24]) );
  CKND2D0 U27 ( .A1(decoder_i[4]), .A2(n7), .ZN(n4) );
  NR2D0 U28 ( .A1(n11), .A2(n5), .ZN(decoder_o[29]) );
  NR2D0 U29 ( .A1(n11), .A2(n14), .ZN(decoder_o[15]) );
  NR2D0 U30 ( .A1(n11), .A2(n16), .ZN(decoder_o[13]) );
  NR2XD0 U31 ( .A1(n3), .A2(n18), .ZN(decoder_o[19]) );
  NR2XD0 U32 ( .A1(n5), .A2(n18), .ZN(decoder_o[17]) );
  ND3D0 U33 ( .A1(decoder_i[1]), .A2(decoder_i[0]), .A3(n9), .ZN(n14) );
  CKND2D1 U34 ( .A1(decoder_i[3]), .A2(n1), .ZN(n12) );
  CKND2D1 U35 ( .A1(decoder_i[2]), .A2(n2), .ZN(n13) );
  CKND2D0 U36 ( .A1(decoder_i[4]), .A2(n10), .ZN(n6) );
  ND3D0 U37 ( .A1(decoder_i[4]), .A2(decoder_i[0]), .A3(n8), .ZN(n5) );
  NR2D0 U38 ( .A1(decoder_i[0]), .A2(n8), .ZN(n7) );
  NR2D0 U39 ( .A1(n11), .A2(n3), .ZN(decoder_o[31]) );
  ND3D0 U40 ( .A1(decoder_i[0]), .A2(n9), .A3(n8), .ZN(n16) );
  CKND0 U41 ( .I(decoder_i[2]), .ZN(n1) );
  ND3D0 U42 ( .A1(decoder_i[4]), .A2(decoder_i[1]), .A3(decoder_i[0]), .ZN(n3)
         );
  NR2D0 U43 ( .A1(decoder_i[1]), .A2(decoder_i[0]), .ZN(n10) );
  CKND2D1 U44 ( .A1(decoder_i[3]), .A2(decoder_i[2]), .ZN(n11) );
  CKND0 U45 ( .I(decoder_i[1]), .ZN(n8) );
  CKND0 U46 ( .I(decoder_i[3]), .ZN(n2) );
  CKND0 U47 ( .I(decoder_i[4]), .ZN(n9) );
  NR2D1 U48 ( .A1(n6), .A2(n18), .ZN(decoder_o[16]) );
  ND2D1 U49 ( .A1(n10), .A2(n9), .ZN(n17) );
  ND2D1 U50 ( .A1(n7), .A2(n9), .ZN(n15) );
endmodule


module priority_encoder ( inp_i, out_o, valid_o );
  input [31:0] inp_i;
  output [4:0] out_o;
  output valid_o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61;

  NR2D1 U1 ( .A1(inp_i[24]), .A2(inp_i[25]), .ZN(n26) );
  NR4D0 U2 ( .A1(inp_i[28]), .A2(inp_i[29]), .A3(inp_i[30]), .A4(inp_i[31]), 
        .ZN(n14) );
  ND2D1 U3 ( .A1(n30), .A2(n26), .ZN(n13) );
  NR2D1 U4 ( .A1(inp_i[18]), .A2(inp_i[19]), .ZN(n27) );
  NR4D0 U5 ( .A1(inp_i[4]), .A2(inp_i[5]), .A3(inp_i[6]), .A4(inp_i[7]), .ZN(
        n19) );
  ND2D1 U6 ( .A1(n25), .A2(n61), .ZN(n15) );
  ND2D1 U7 ( .A1(n60), .A2(n24), .ZN(n18) );
  NR2D1 U8 ( .A1(inp_i[10]), .A2(inp_i[11]), .ZN(n60) );
  NR2D1 U9 ( .A1(inp_i[14]), .A2(inp_i[15]), .ZN(n61) );
  INVD1 U10 ( .I(n13), .ZN(n10) );
  INR2D1 U11 ( .A1(n19), .B1(n17), .ZN(n11) );
  IND3D1 U12 ( .A1(n9), .B1(n10), .B2(n14), .ZN(n59) );
  AOI221D1 U13 ( .A1(inp_i[6]), .A2(n55), .B1(n54), .B2(n55), .C(inp_i[0]), 
        .ZN(out_o[0]) );
  AOI221D0 U14 ( .A1(inp_i[3]), .A2(n43), .B1(n42), .B2(n43), .C(inp_i[1]), 
        .ZN(n55) );
  AOI221D1 U15 ( .A1(inp_i[1]), .A2(n39), .B1(n38), .B2(n39), .C(inp_i[0]), 
        .ZN(out_o[1]) );
  AOI32D1 U16 ( .A1(n34), .A2(n57), .A3(n56), .B1(n33), .B2(n57), .ZN(n39) );
  AOI221D1 U17 ( .A1(n20), .A2(n19), .B1(n18), .B2(n19), .C(n17), .ZN(out_o[2]) );
  AOI221D0 U18 ( .A1(inp_i[25]), .A2(n47), .B1(n46), .B2(n47), .C(inp_i[23]), 
        .ZN(n1) );
  AOI221D0 U19 ( .A1(n1), .A2(n48), .B1(inp_i[22]), .B2(n48), .C(inp_i[20]), 
        .ZN(n49) );
  CKND0 U20 ( .I(inp_i[13]), .ZN(n2) );
  AOI221D0 U21 ( .A1(inp_i[14]), .A2(n2), .B1(n51), .B2(n2), .C(inp_i[12]), 
        .ZN(n52) );
  AOI211D0 U22 ( .A1(n10), .A2(n14), .B(inp_i[16]), .C(n9), .ZN(n3) );
  OA31D0 U23 ( .A1(n3), .A2(n15), .A3(n18), .B(n11), .Z(out_o[3]) );
  AOI21D0 U24 ( .A1(inp_i[31]), .A2(n44), .B(inp_i[29]), .ZN(n4) );
  AOI221D0 U25 ( .A1(inp_i[28]), .A2(n45), .B1(n4), .B2(n45), .C(inp_i[26]), 
        .ZN(n46) );
  OAI21D0 U26 ( .A1(n59), .A2(inp_i[16]), .B(n11), .ZN(n5) );
  NR3D0 U27 ( .A1(n15), .A2(n18), .A3(n5), .ZN(out_o[4]) );
  CKND0 U28 ( .I(inp_i[10]), .ZN(n6) );
  AOI221D0 U29 ( .A1(inp_i[11]), .A2(n6), .B1(n52), .B2(n6), .C(inp_i[9]), 
        .ZN(n53) );
  ND3D0 U30 ( .A1(n56), .A2(n57), .A3(n58), .ZN(n7) );
  NR4D0 U31 ( .A1(n59), .A2(inp_i[2]), .A3(inp_i[3]), .A4(n7), .ZN(n8) );
  IND4D0 U32 ( .A1(inp_i[0]), .B1(n60), .B2(n8), .B3(n61), .ZN(valid_o) );
  OR4D1 U33 ( .A1(inp_i[2]), .A2(inp_i[4]), .A3(n53), .A4(inp_i[8]), .Z(n54)
         );
  IAO21D0 U34 ( .A1(inp_i[19]), .A2(n49), .B(inp_i[18]), .ZN(n50) );
  AOI211XD0 U35 ( .A1(n37), .A2(n36), .B(inp_i[2]), .C(inp_i[3]), .ZN(n38) );
  OAI21D0 U36 ( .A1(n60), .A2(n35), .B(n58), .ZN(n36) );
  OAI21D0 U37 ( .A1(n14), .A2(n13), .B(n12), .ZN(n16) );
  AOI211XD0 U38 ( .A1(n23), .A2(n22), .B(inp_i[17]), .C(n28), .ZN(n34) );
  NR2D0 U39 ( .A1(inp_i[4]), .A2(n41), .ZN(n42) );
  INVD0 U40 ( .I(n24), .ZN(n35) );
  AOI21D0 U41 ( .A1(inp_i[7]), .A2(n40), .B(inp_i[5]), .ZN(n41) );
  OAI211D0 U42 ( .A1(inp_i[30]), .A2(inp_i[31]), .B(n26), .C(n21), .ZN(n22) );
  CKND0 U43 ( .I(n26), .ZN(n29) );
  CKND1 U44 ( .I(inp_i[2]), .ZN(n43) );
  NR2D0 U45 ( .A1(inp_i[6]), .A2(inp_i[7]), .ZN(n58) );
  NR2D0 U46 ( .A1(inp_i[16]), .A2(inp_i[17]), .ZN(n32) );
  OR4D1 U47 ( .A1(inp_i[0]), .A2(inp_i[1]), .A3(inp_i[2]), .A4(inp_i[3]), .Z(
        n17) );
  NR2D0 U48 ( .A1(inp_i[22]), .A2(inp_i[23]), .ZN(n23) );
  CKND1 U49 ( .I(inp_i[21]), .ZN(n48) );
  NR2D0 U50 ( .A1(inp_i[28]), .A2(inp_i[29]), .ZN(n21) );
  NR2D0 U51 ( .A1(inp_i[4]), .A2(inp_i[5]), .ZN(n37) );
  CKND0 U52 ( .I(inp_i[30]), .ZN(n44) );
  CKND0 U53 ( .I(inp_i[27]), .ZN(n45) );
  CKND0 U54 ( .I(inp_i[24]), .ZN(n47) );
  CKND0 U55 ( .I(inp_i[6]), .ZN(n40) );
  AOI31D1 U56 ( .A1(n27), .A2(n32), .A3(n16), .B(n15), .ZN(n20) );
  NR2D1 U57 ( .A1(inp_i[26]), .A2(inp_i[27]), .ZN(n30) );
  NR2D1 U58 ( .A1(inp_i[9]), .A2(inp_i[8]), .ZN(n24) );
  NR2D1 U59 ( .A1(inp_i[12]), .A2(inp_i[13]), .ZN(n25) );
  INVD1 U60 ( .I(inp_i[16]), .ZN(n56) );
  IND3D1 U61 ( .A1(inp_i[17]), .B1(n27), .B2(n12), .ZN(n9) );
  IOA21D1 U62 ( .A1(n32), .A2(n31), .B(n61), .ZN(n33) );
  OAI31D1 U63 ( .A1(n30), .A2(n29), .A3(n28), .B(n27), .ZN(n31) );
  IND2D1 U64 ( .A1(inp_i[20]), .B1(n48), .ZN(n28) );
  NR4D0 U65 ( .A1(inp_i[20]), .A2(inp_i[21]), .A3(inp_i[22]), .A4(inp_i[23]), 
        .ZN(n12) );
  IINR4D0 U66 ( .A1(n25), .A2(n37), .B1(n35), .B2(inp_i[1]), .ZN(n57) );
  AOI221D0 U67 ( .A1(inp_i[17]), .A2(n56), .B1(n50), .B2(n56), .C(inp_i[15]), 
        .ZN(n51) );
endmodule


module mux ( .data_i({\data_i[31][31] , \data_i[31][30] , \data_i[31][29] , 
        \data_i[31][28] , \data_i[31][27] , \data_i[31][26] , \data_i[31][25] , 
        \data_i[31][24] , \data_i[31][23] , \data_i[31][22] , \data_i[31][21] , 
        \data_i[31][20] , \data_i[31][19] , \data_i[31][18] , \data_i[31][17] , 
        \data_i[31][16] , \data_i[31][15] , \data_i[31][14] , \data_i[31][13] , 
        \data_i[31][12] , \data_i[31][11] , \data_i[31][10] , \data_i[31][9] , 
        \data_i[31][8] , \data_i[31][7] , \data_i[31][6] , \data_i[31][5] , 
        \data_i[31][4] , \data_i[31][3] , \data_i[31][2] , \data_i[31][1] , 
        \data_i[31][0] , \data_i[30][31] , \data_i[30][30] , \data_i[30][29] , 
        \data_i[30][28] , \data_i[30][27] , \data_i[30][26] , \data_i[30][25] , 
        \data_i[30][24] , \data_i[30][23] , \data_i[30][22] , \data_i[30][21] , 
        \data_i[30][20] , \data_i[30][19] , \data_i[30][18] , \data_i[30][17] , 
        \data_i[30][16] , \data_i[30][15] , \data_i[30][14] , \data_i[30][13] , 
        \data_i[30][12] , \data_i[30][11] , \data_i[30][10] , \data_i[30][9] , 
        \data_i[30][8] , \data_i[30][7] , \data_i[30][6] , \data_i[30][5] , 
        \data_i[30][4] , \data_i[30][3] , \data_i[30][2] , \data_i[30][1] , 
        \data_i[30][0] , \data_i[29][31] , \data_i[29][30] , \data_i[29][29] , 
        \data_i[29][28] , \data_i[29][27] , \data_i[29][26] , \data_i[29][25] , 
        \data_i[29][24] , \data_i[29][23] , \data_i[29][22] , \data_i[29][21] , 
        \data_i[29][20] , \data_i[29][19] , \data_i[29][18] , \data_i[29][17] , 
        \data_i[29][16] , \data_i[29][15] , \data_i[29][14] , \data_i[29][13] , 
        \data_i[29][12] , \data_i[29][11] , \data_i[29][10] , \data_i[29][9] , 
        \data_i[29][8] , \data_i[29][7] , \data_i[29][6] , \data_i[29][5] , 
        \data_i[29][4] , \data_i[29][3] , \data_i[29][2] , \data_i[29][1] , 
        \data_i[29][0] , \data_i[28][31] , \data_i[28][30] , \data_i[28][29] , 
        \data_i[28][28] , \data_i[28][27] , \data_i[28][26] , \data_i[28][25] , 
        \data_i[28][24] , \data_i[28][23] , \data_i[28][22] , \data_i[28][21] , 
        \data_i[28][20] , \data_i[28][19] , \data_i[28][18] , \data_i[28][17] , 
        \data_i[28][16] , \data_i[28][15] , \data_i[28][14] , \data_i[28][13] , 
        \data_i[28][12] , \data_i[28][11] , \data_i[28][10] , \data_i[28][9] , 
        \data_i[28][8] , \data_i[28][7] , \data_i[28][6] , \data_i[28][5] , 
        \data_i[28][4] , \data_i[28][3] , \data_i[28][2] , \data_i[28][1] , 
        \data_i[28][0] , \data_i[27][31] , \data_i[27][30] , \data_i[27][29] , 
        \data_i[27][28] , \data_i[27][27] , \data_i[27][26] , \data_i[27][25] , 
        \data_i[27][24] , \data_i[27][23] , \data_i[27][22] , \data_i[27][21] , 
        \data_i[27][20] , \data_i[27][19] , \data_i[27][18] , \data_i[27][17] , 
        \data_i[27][16] , \data_i[27][15] , \data_i[27][14] , \data_i[27][13] , 
        \data_i[27][12] , \data_i[27][11] , \data_i[27][10] , \data_i[27][9] , 
        \data_i[27][8] , \data_i[27][7] , \data_i[27][6] , \data_i[27][5] , 
        \data_i[27][4] , \data_i[27][3] , \data_i[27][2] , \data_i[27][1] , 
        \data_i[27][0] , \data_i[26][31] , \data_i[26][30] , \data_i[26][29] , 
        \data_i[26][28] , \data_i[26][27] , \data_i[26][26] , \data_i[26][25] , 
        \data_i[26][24] , \data_i[26][23] , \data_i[26][22] , \data_i[26][21] , 
        \data_i[26][20] , \data_i[26][19] , \data_i[26][18] , \data_i[26][17] , 
        \data_i[26][16] , \data_i[26][15] , \data_i[26][14] , \data_i[26][13] , 
        \data_i[26][12] , \data_i[26][11] , \data_i[26][10] , \data_i[26][9] , 
        \data_i[26][8] , \data_i[26][7] , \data_i[26][6] , \data_i[26][5] , 
        \data_i[26][4] , \data_i[26][3] , \data_i[26][2] , \data_i[26][1] , 
        \data_i[26][0] , \data_i[25][31] , \data_i[25][30] , \data_i[25][29] , 
        \data_i[25][28] , \data_i[25][27] , \data_i[25][26] , \data_i[25][25] , 
        \data_i[25][24] , \data_i[25][23] , \data_i[25][22] , \data_i[25][21] , 
        \data_i[25][20] , \data_i[25][19] , \data_i[25][18] , \data_i[25][17] , 
        \data_i[25][16] , \data_i[25][15] , \data_i[25][14] , \data_i[25][13] , 
        \data_i[25][12] , \data_i[25][11] , \data_i[25][10] , \data_i[25][9] , 
        \data_i[25][8] , \data_i[25][7] , \data_i[25][6] , \data_i[25][5] , 
        \data_i[25][4] , \data_i[25][3] , \data_i[25][2] , \data_i[25][1] , 
        \data_i[25][0] , \data_i[24][31] , \data_i[24][30] , \data_i[24][29] , 
        \data_i[24][28] , \data_i[24][27] , \data_i[24][26] , \data_i[24][25] , 
        \data_i[24][24] , \data_i[24][23] , \data_i[24][22] , \data_i[24][21] , 
        \data_i[24][20] , \data_i[24][19] , \data_i[24][18] , \data_i[24][17] , 
        \data_i[24][16] , \data_i[24][15] , \data_i[24][14] , \data_i[24][13] , 
        \data_i[24][12] , \data_i[24][11] , \data_i[24][10] , \data_i[24][9] , 
        \data_i[24][8] , \data_i[24][7] , \data_i[24][6] , \data_i[24][5] , 
        \data_i[24][4] , \data_i[24][3] , \data_i[24][2] , \data_i[24][1] , 
        \data_i[24][0] , \data_i[23][31] , \data_i[23][30] , \data_i[23][29] , 
        \data_i[23][28] , \data_i[23][27] , \data_i[23][26] , \data_i[23][25] , 
        \data_i[23][24] , \data_i[23][23] , \data_i[23][22] , \data_i[23][21] , 
        \data_i[23][20] , \data_i[23][19] , \data_i[23][18] , \data_i[23][17] , 
        \data_i[23][16] , \data_i[23][15] , \data_i[23][14] , \data_i[23][13] , 
        \data_i[23][12] , \data_i[23][11] , \data_i[23][10] , \data_i[23][9] , 
        \data_i[23][8] , \data_i[23][7] , \data_i[23][6] , \data_i[23][5] , 
        \data_i[23][4] , \data_i[23][3] , \data_i[23][2] , \data_i[23][1] , 
        \data_i[23][0] , \data_i[22][31] , \data_i[22][30] , \data_i[22][29] , 
        \data_i[22][28] , \data_i[22][27] , \data_i[22][26] , \data_i[22][25] , 
        \data_i[22][24] , \data_i[22][23] , \data_i[22][22] , \data_i[22][21] , 
        \data_i[22][20] , \data_i[22][19] , \data_i[22][18] , \data_i[22][17] , 
        \data_i[22][16] , \data_i[22][15] , \data_i[22][14] , \data_i[22][13] , 
        \data_i[22][12] , \data_i[22][11] , \data_i[22][10] , \data_i[22][9] , 
        \data_i[22][8] , \data_i[22][7] , \data_i[22][6] , \data_i[22][5] , 
        \data_i[22][4] , \data_i[22][3] , \data_i[22][2] , \data_i[22][1] , 
        \data_i[22][0] , \data_i[21][31] , \data_i[21][30] , \data_i[21][29] , 
        \data_i[21][28] , \data_i[21][27] , \data_i[21][26] , \data_i[21][25] , 
        \data_i[21][24] , \data_i[21][23] , \data_i[21][22] , \data_i[21][21] , 
        \data_i[21][20] , \data_i[21][19] , \data_i[21][18] , \data_i[21][17] , 
        \data_i[21][16] , \data_i[21][15] , \data_i[21][14] , \data_i[21][13] , 
        \data_i[21][12] , \data_i[21][11] , \data_i[21][10] , \data_i[21][9] , 
        \data_i[21][8] , \data_i[21][7] , \data_i[21][6] , \data_i[21][5] , 
        \data_i[21][4] , \data_i[21][3] , \data_i[21][2] , \data_i[21][1] , 
        \data_i[21][0] , \data_i[20][31] , \data_i[20][30] , \data_i[20][29] , 
        \data_i[20][28] , \data_i[20][27] , \data_i[20][26] , \data_i[20][25] , 
        \data_i[20][24] , \data_i[20][23] , \data_i[20][22] , \data_i[20][21] , 
        \data_i[20][20] , \data_i[20][19] , \data_i[20][18] , \data_i[20][17] , 
        \data_i[20][16] , \data_i[20][15] , \data_i[20][14] , \data_i[20][13] , 
        \data_i[20][12] , \data_i[20][11] , \data_i[20][10] , \data_i[20][9] , 
        \data_i[20][8] , \data_i[20][7] , \data_i[20][6] , \data_i[20][5] , 
        \data_i[20][4] , \data_i[20][3] , \data_i[20][2] , \data_i[20][1] , 
        \data_i[20][0] , \data_i[19][31] , \data_i[19][30] , \data_i[19][29] , 
        \data_i[19][28] , \data_i[19][27] , \data_i[19][26] , \data_i[19][25] , 
        \data_i[19][24] , \data_i[19][23] , \data_i[19][22] , \data_i[19][21] , 
        \data_i[19][20] , \data_i[19][19] , \data_i[19][18] , \data_i[19][17] , 
        \data_i[19][16] , \data_i[19][15] , \data_i[19][14] , \data_i[19][13] , 
        \data_i[19][12] , \data_i[19][11] , \data_i[19][10] , \data_i[19][9] , 
        \data_i[19][8] , \data_i[19][7] , \data_i[19][6] , \data_i[19][5] , 
        \data_i[19][4] , \data_i[19][3] , \data_i[19][2] , \data_i[19][1] , 
        \data_i[19][0] , \data_i[18][31] , \data_i[18][30] , \data_i[18][29] , 
        \data_i[18][28] , \data_i[18][27] , \data_i[18][26] , \data_i[18][25] , 
        \data_i[18][24] , \data_i[18][23] , \data_i[18][22] , \data_i[18][21] , 
        \data_i[18][20] , \data_i[18][19] , \data_i[18][18] , \data_i[18][17] , 
        \data_i[18][16] , \data_i[18][15] , \data_i[18][14] , \data_i[18][13] , 
        \data_i[18][12] , \data_i[18][11] , \data_i[18][10] , \data_i[18][9] , 
        \data_i[18][8] , \data_i[18][7] , \data_i[18][6] , \data_i[18][5] , 
        \data_i[18][4] , \data_i[18][3] , \data_i[18][2] , \data_i[18][1] , 
        \data_i[18][0] , \data_i[17][31] , \data_i[17][30] , \data_i[17][29] , 
        \data_i[17][28] , \data_i[17][27] , \data_i[17][26] , \data_i[17][25] , 
        \data_i[17][24] , \data_i[17][23] , \data_i[17][22] , \data_i[17][21] , 
        \data_i[17][20] , \data_i[17][19] , \data_i[17][18] , \data_i[17][17] , 
        \data_i[17][16] , \data_i[17][15] , \data_i[17][14] , \data_i[17][13] , 
        \data_i[17][12] , \data_i[17][11] , \data_i[17][10] , \data_i[17][9] , 
        \data_i[17][8] , \data_i[17][7] , \data_i[17][6] , \data_i[17][5] , 
        \data_i[17][4] , \data_i[17][3] , \data_i[17][2] , \data_i[17][1] , 
        \data_i[17][0] , \data_i[16][31] , \data_i[16][30] , \data_i[16][29] , 
        \data_i[16][28] , \data_i[16][27] , \data_i[16][26] , \data_i[16][25] , 
        \data_i[16][24] , \data_i[16][23] , \data_i[16][22] , \data_i[16][21] , 
        \data_i[16][20] , \data_i[16][19] , \data_i[16][18] , \data_i[16][17] , 
        \data_i[16][16] , \data_i[16][15] , \data_i[16][14] , \data_i[16][13] , 
        \data_i[16][12] , \data_i[16][11] , \data_i[16][10] , \data_i[16][9] , 
        \data_i[16][8] , \data_i[16][7] , \data_i[16][6] , \data_i[16][5] , 
        \data_i[16][4] , \data_i[16][3] , \data_i[16][2] , \data_i[16][1] , 
        \data_i[16][0] , \data_i[15][31] , \data_i[15][30] , \data_i[15][29] , 
        \data_i[15][28] , \data_i[15][27] , \data_i[15][26] , \data_i[15][25] , 
        \data_i[15][24] , \data_i[15][23] , \data_i[15][22] , \data_i[15][21] , 
        \data_i[15][20] , \data_i[15][19] , \data_i[15][18] , \data_i[15][17] , 
        \data_i[15][16] , \data_i[15][15] , \data_i[15][14] , \data_i[15][13] , 
        \data_i[15][12] , \data_i[15][11] , \data_i[15][10] , \data_i[15][9] , 
        \data_i[15][8] , \data_i[15][7] , \data_i[15][6] , \data_i[15][5] , 
        \data_i[15][4] , \data_i[15][3] , \data_i[15][2] , \data_i[15][1] , 
        \data_i[15][0] , \data_i[14][31] , \data_i[14][30] , \data_i[14][29] , 
        \data_i[14][28] , \data_i[14][27] , \data_i[14][26] , \data_i[14][25] , 
        \data_i[14][24] , \data_i[14][23] , \data_i[14][22] , \data_i[14][21] , 
        \data_i[14][20] , \data_i[14][19] , \data_i[14][18] , \data_i[14][17] , 
        \data_i[14][16] , \data_i[14][15] , \data_i[14][14] , \data_i[14][13] , 
        \data_i[14][12] , \data_i[14][11] , \data_i[14][10] , \data_i[14][9] , 
        \data_i[14][8] , \data_i[14][7] , \data_i[14][6] , \data_i[14][5] , 
        \data_i[14][4] , \data_i[14][3] , \data_i[14][2] , \data_i[14][1] , 
        \data_i[14][0] , \data_i[13][31] , \data_i[13][30] , \data_i[13][29] , 
        \data_i[13][28] , \data_i[13][27] , \data_i[13][26] , \data_i[13][25] , 
        \data_i[13][24] , \data_i[13][23] , \data_i[13][22] , \data_i[13][21] , 
        \data_i[13][20] , \data_i[13][19] , \data_i[13][18] , \data_i[13][17] , 
        \data_i[13][16] , \data_i[13][15] , \data_i[13][14] , \data_i[13][13] , 
        \data_i[13][12] , \data_i[13][11] , \data_i[13][10] , \data_i[13][9] , 
        \data_i[13][8] , \data_i[13][7] , \data_i[13][6] , \data_i[13][5] , 
        \data_i[13][4] , \data_i[13][3] , \data_i[13][2] , \data_i[13][1] , 
        \data_i[13][0] , \data_i[12][31] , \data_i[12][30] , \data_i[12][29] , 
        \data_i[12][28] , \data_i[12][27] , \data_i[12][26] , \data_i[12][25] , 
        \data_i[12][24] , \data_i[12][23] , \data_i[12][22] , \data_i[12][21] , 
        \data_i[12][20] , \data_i[12][19] , \data_i[12][18] , \data_i[12][17] , 
        \data_i[12][16] , \data_i[12][15] , \data_i[12][14] , \data_i[12][13] , 
        \data_i[12][12] , \data_i[12][11] , \data_i[12][10] , \data_i[12][9] , 
        \data_i[12][8] , \data_i[12][7] , \data_i[12][6] , \data_i[12][5] , 
        \data_i[12][4] , \data_i[12][3] , \data_i[12][2] , \data_i[12][1] , 
        \data_i[12][0] , \data_i[11][31] , \data_i[11][30] , \data_i[11][29] , 
        \data_i[11][28] , \data_i[11][27] , \data_i[11][26] , \data_i[11][25] , 
        \data_i[11][24] , \data_i[11][23] , \data_i[11][22] , \data_i[11][21] , 
        \data_i[11][20] , \data_i[11][19] , \data_i[11][18] , \data_i[11][17] , 
        \data_i[11][16] , \data_i[11][15] , \data_i[11][14] , \data_i[11][13] , 
        \data_i[11][12] , \data_i[11][11] , \data_i[11][10] , \data_i[11][9] , 
        \data_i[11][8] , \data_i[11][7] , \data_i[11][6] , \data_i[11][5] , 
        \data_i[11][4] , \data_i[11][3] , \data_i[11][2] , \data_i[11][1] , 
        \data_i[11][0] , \data_i[10][31] , \data_i[10][30] , \data_i[10][29] , 
        \data_i[10][28] , \data_i[10][27] , \data_i[10][26] , \data_i[10][25] , 
        \data_i[10][24] , \data_i[10][23] , \data_i[10][22] , \data_i[10][21] , 
        \data_i[10][20] , \data_i[10][19] , \data_i[10][18] , \data_i[10][17] , 
        \data_i[10][16] , \data_i[10][15] , \data_i[10][14] , \data_i[10][13] , 
        \data_i[10][12] , \data_i[10][11] , \data_i[10][10] , \data_i[10][9] , 
        \data_i[10][8] , \data_i[10][7] , \data_i[10][6] , \data_i[10][5] , 
        \data_i[10][4] , \data_i[10][3] , \data_i[10][2] , \data_i[10][1] , 
        \data_i[10][0] , \data_i[9][31] , \data_i[9][30] , \data_i[9][29] , 
        \data_i[9][28] , \data_i[9][27] , \data_i[9][26] , \data_i[9][25] , 
        \data_i[9][24] , \data_i[9][23] , \data_i[9][22] , \data_i[9][21] , 
        \data_i[9][20] , \data_i[9][19] , \data_i[9][18] , \data_i[9][17] , 
        \data_i[9][16] , \data_i[9][15] , \data_i[9][14] , \data_i[9][13] , 
        \data_i[9][12] , \data_i[9][11] , \data_i[9][10] , \data_i[9][9] , 
        \data_i[9][8] , \data_i[9][7] , \data_i[9][6] , \data_i[9][5] , 
        \data_i[9][4] , \data_i[9][3] , \data_i[9][2] , \data_i[9][1] , 
        \data_i[9][0] , \data_i[8][31] , \data_i[8][30] , \data_i[8][29] , 
        \data_i[8][28] , \data_i[8][27] , \data_i[8][26] , \data_i[8][25] , 
        \data_i[8][24] , \data_i[8][23] , \data_i[8][22] , \data_i[8][21] , 
        \data_i[8][20] , \data_i[8][19] , \data_i[8][18] , \data_i[8][17] , 
        \data_i[8][16] , \data_i[8][15] , \data_i[8][14] , \data_i[8][13] , 
        \data_i[8][12] , \data_i[8][11] , \data_i[8][10] , \data_i[8][9] , 
        \data_i[8][8] , \data_i[8][7] , \data_i[8][6] , \data_i[8][5] , 
        \data_i[8][4] , \data_i[8][3] , \data_i[8][2] , \data_i[8][1] , 
        \data_i[8][0] , \data_i[7][31] , \data_i[7][30] , \data_i[7][29] , 
        \data_i[7][28] , \data_i[7][27] , \data_i[7][26] , \data_i[7][25] , 
        \data_i[7][24] , \data_i[7][23] , \data_i[7][22] , \data_i[7][21] , 
        \data_i[7][20] , \data_i[7][19] , \data_i[7][18] , \data_i[7][17] , 
        \data_i[7][16] , \data_i[7][15] , \data_i[7][14] , \data_i[7][13] , 
        \data_i[7][12] , \data_i[7][11] , \data_i[7][10] , \data_i[7][9] , 
        \data_i[7][8] , \data_i[7][7] , \data_i[7][6] , \data_i[7][5] , 
        \data_i[7][4] , \data_i[7][3] , \data_i[7][2] , \data_i[7][1] , 
        \data_i[7][0] , \data_i[6][31] , \data_i[6][30] , \data_i[6][29] , 
        \data_i[6][28] , \data_i[6][27] , \data_i[6][26] , \data_i[6][25] , 
        \data_i[6][24] , \data_i[6][23] , \data_i[6][22] , \data_i[6][21] , 
        \data_i[6][20] , \data_i[6][19] , \data_i[6][18] , \data_i[6][17] , 
        \data_i[6][16] , \data_i[6][15] , \data_i[6][14] , \data_i[6][13] , 
        \data_i[6][12] , \data_i[6][11] , \data_i[6][10] , \data_i[6][9] , 
        \data_i[6][8] , \data_i[6][7] , \data_i[6][6] , \data_i[6][5] , 
        \data_i[6][4] , \data_i[6][3] , \data_i[6][2] , \data_i[6][1] , 
        \data_i[6][0] , \data_i[5][31] , \data_i[5][30] , \data_i[5][29] , 
        \data_i[5][28] , \data_i[5][27] , \data_i[5][26] , \data_i[5][25] , 
        \data_i[5][24] , \data_i[5][23] , \data_i[5][22] , \data_i[5][21] , 
        \data_i[5][20] , \data_i[5][19] , \data_i[5][18] , \data_i[5][17] , 
        \data_i[5][16] , \data_i[5][15] , \data_i[5][14] , \data_i[5][13] , 
        \data_i[5][12] , \data_i[5][11] , \data_i[5][10] , \data_i[5][9] , 
        \data_i[5][8] , \data_i[5][7] , \data_i[5][6] , \data_i[5][5] , 
        \data_i[5][4] , \data_i[5][3] , \data_i[5][2] , \data_i[5][1] , 
        \data_i[5][0] , \data_i[4][31] , \data_i[4][30] , \data_i[4][29] , 
        \data_i[4][28] , \data_i[4][27] , \data_i[4][26] , \data_i[4][25] , 
        \data_i[4][24] , \data_i[4][23] , \data_i[4][22] , \data_i[4][21] , 
        \data_i[4][20] , \data_i[4][19] , \data_i[4][18] , \data_i[4][17] , 
        \data_i[4][16] , \data_i[4][15] , \data_i[4][14] , \data_i[4][13] , 
        \data_i[4][12] , \data_i[4][11] , \data_i[4][10] , \data_i[4][9] , 
        \data_i[4][8] , \data_i[4][7] , \data_i[4][6] , \data_i[4][5] , 
        \data_i[4][4] , \data_i[4][3] , \data_i[4][2] , \data_i[4][1] , 
        \data_i[4][0] , \data_i[3][31] , \data_i[3][30] , \data_i[3][29] , 
        \data_i[3][28] , \data_i[3][27] , \data_i[3][26] , \data_i[3][25] , 
        \data_i[3][24] , \data_i[3][23] , \data_i[3][22] , \data_i[3][21] , 
        \data_i[3][20] , \data_i[3][19] , \data_i[3][18] , \data_i[3][17] , 
        \data_i[3][16] , \data_i[3][15] , \data_i[3][14] , \data_i[3][13] , 
        \data_i[3][12] , \data_i[3][11] , \data_i[3][10] , \data_i[3][9] , 
        \data_i[3][8] , \data_i[3][7] , \data_i[3][6] , \data_i[3][5] , 
        \data_i[3][4] , \data_i[3][3] , \data_i[3][2] , \data_i[3][1] , 
        \data_i[3][0] , \data_i[2][31] , \data_i[2][30] , \data_i[2][29] , 
        \data_i[2][28] , \data_i[2][27] , \data_i[2][26] , \data_i[2][25] , 
        \data_i[2][24] , \data_i[2][23] , \data_i[2][22] , \data_i[2][21] , 
        \data_i[2][20] , \data_i[2][19] , \data_i[2][18] , \data_i[2][17] , 
        \data_i[2][16] , \data_i[2][15] , \data_i[2][14] , \data_i[2][13] , 
        \data_i[2][12] , \data_i[2][11] , \data_i[2][10] , \data_i[2][9] , 
        \data_i[2][8] , \data_i[2][7] , \data_i[2][6] , \data_i[2][5] , 
        \data_i[2][4] , \data_i[2][3] , \data_i[2][2] , \data_i[2][1] , 
        \data_i[2][0] , \data_i[1][31] , \data_i[1][30] , \data_i[1][29] , 
        \data_i[1][28] , \data_i[1][27] , \data_i[1][26] , \data_i[1][25] , 
        \data_i[1][24] , \data_i[1][23] , \data_i[1][22] , \data_i[1][21] , 
        \data_i[1][20] , \data_i[1][19] , \data_i[1][18] , \data_i[1][17] , 
        \data_i[1][16] , \data_i[1][15] , \data_i[1][14] , \data_i[1][13] , 
        \data_i[1][12] , \data_i[1][11] , \data_i[1][10] , \data_i[1][9] , 
        \data_i[1][8] , \data_i[1][7] , \data_i[1][6] , \data_i[1][5] , 
        \data_i[1][4] , \data_i[1][3] , \data_i[1][2] , \data_i[1][1] , 
        \data_i[1][0] , \data_i[0][31] , \data_i[0][30] , \data_i[0][29] , 
        \data_i[0][28] , \data_i[0][27] , \data_i[0][26] , \data_i[0][25] , 
        \data_i[0][24] , \data_i[0][23] , \data_i[0][22] , \data_i[0][21] , 
        \data_i[0][20] , \data_i[0][19] , \data_i[0][18] , \data_i[0][17] , 
        \data_i[0][16] , \data_i[0][15] , \data_i[0][14] , \data_i[0][13] , 
        \data_i[0][12] , \data_i[0][11] , \data_i[0][10] , \data_i[0][9] , 
        \data_i[0][8] , \data_i[0][7] , \data_i[0][6] , \data_i[0][5] , 
        \data_i[0][4] , \data_i[0][3] , \data_i[0][2] , \data_i[0][1] , 
        \data_i[0][0] }), select_i, data_o );
  input [4:0] select_i;
  output [31:0] data_o;
  input \data_i[31][31] , \data_i[31][30] , \data_i[31][29] , \data_i[31][28] ,
         \data_i[31][27] , \data_i[31][26] , \data_i[31][25] ,
         \data_i[31][24] , \data_i[31][23] , \data_i[31][22] ,
         \data_i[31][21] , \data_i[31][20] , \data_i[31][19] ,
         \data_i[31][18] , \data_i[31][17] , \data_i[31][16] ,
         \data_i[31][15] , \data_i[31][14] , \data_i[31][13] ,
         \data_i[31][12] , \data_i[31][11] , \data_i[31][10] , \data_i[31][9] ,
         \data_i[31][8] , \data_i[31][7] , \data_i[31][6] , \data_i[31][5] ,
         \data_i[31][4] , \data_i[31][3] , \data_i[31][2] , \data_i[31][1] ,
         \data_i[31][0] , \data_i[30][31] , \data_i[30][30] , \data_i[30][29] ,
         \data_i[30][28] , \data_i[30][27] , \data_i[30][26] ,
         \data_i[30][25] , \data_i[30][24] , \data_i[30][23] ,
         \data_i[30][22] , \data_i[30][21] , \data_i[30][20] ,
         \data_i[30][19] , \data_i[30][18] , \data_i[30][17] ,
         \data_i[30][16] , \data_i[30][15] , \data_i[30][14] ,
         \data_i[30][13] , \data_i[30][12] , \data_i[30][11] ,
         \data_i[30][10] , \data_i[30][9] , \data_i[30][8] , \data_i[30][7] ,
         \data_i[30][6] , \data_i[30][5] , \data_i[30][4] , \data_i[30][3] ,
         \data_i[30][2] , \data_i[30][1] , \data_i[30][0] , \data_i[29][31] ,
         \data_i[29][30] , \data_i[29][29] , \data_i[29][28] ,
         \data_i[29][27] , \data_i[29][26] , \data_i[29][25] ,
         \data_i[29][24] , \data_i[29][23] , \data_i[29][22] ,
         \data_i[29][21] , \data_i[29][20] , \data_i[29][19] ,
         \data_i[29][18] , \data_i[29][17] , \data_i[29][16] ,
         \data_i[29][15] , \data_i[29][14] , \data_i[29][13] ,
         \data_i[29][12] , \data_i[29][11] , \data_i[29][10] , \data_i[29][9] ,
         \data_i[29][8] , \data_i[29][7] , \data_i[29][6] , \data_i[29][5] ,
         \data_i[29][4] , \data_i[29][3] , \data_i[29][2] , \data_i[29][1] ,
         \data_i[29][0] , \data_i[28][31] , \data_i[28][30] , \data_i[28][29] ,
         \data_i[28][28] , \data_i[28][27] , \data_i[28][26] ,
         \data_i[28][25] , \data_i[28][24] , \data_i[28][23] ,
         \data_i[28][22] , \data_i[28][21] , \data_i[28][20] ,
         \data_i[28][19] , \data_i[28][18] , \data_i[28][17] ,
         \data_i[28][16] , \data_i[28][15] , \data_i[28][14] ,
         \data_i[28][13] , \data_i[28][12] , \data_i[28][11] ,
         \data_i[28][10] , \data_i[28][9] , \data_i[28][8] , \data_i[28][7] ,
         \data_i[28][6] , \data_i[28][5] , \data_i[28][4] , \data_i[28][3] ,
         \data_i[28][2] , \data_i[28][1] , \data_i[28][0] , \data_i[27][31] ,
         \data_i[27][30] , \data_i[27][29] , \data_i[27][28] ,
         \data_i[27][27] , \data_i[27][26] , \data_i[27][25] ,
         \data_i[27][24] , \data_i[27][23] , \data_i[27][22] ,
         \data_i[27][21] , \data_i[27][20] , \data_i[27][19] ,
         \data_i[27][18] , \data_i[27][17] , \data_i[27][16] ,
         \data_i[27][15] , \data_i[27][14] , \data_i[27][13] ,
         \data_i[27][12] , \data_i[27][11] , \data_i[27][10] , \data_i[27][9] ,
         \data_i[27][8] , \data_i[27][7] , \data_i[27][6] , \data_i[27][5] ,
         \data_i[27][4] , \data_i[27][3] , \data_i[27][2] , \data_i[27][1] ,
         \data_i[27][0] , \data_i[26][31] , \data_i[26][30] , \data_i[26][29] ,
         \data_i[26][28] , \data_i[26][27] , \data_i[26][26] ,
         \data_i[26][25] , \data_i[26][24] , \data_i[26][23] ,
         \data_i[26][22] , \data_i[26][21] , \data_i[26][20] ,
         \data_i[26][19] , \data_i[26][18] , \data_i[26][17] ,
         \data_i[26][16] , \data_i[26][15] , \data_i[26][14] ,
         \data_i[26][13] , \data_i[26][12] , \data_i[26][11] ,
         \data_i[26][10] , \data_i[26][9] , \data_i[26][8] , \data_i[26][7] ,
         \data_i[26][6] , \data_i[26][5] , \data_i[26][4] , \data_i[26][3] ,
         \data_i[26][2] , \data_i[26][1] , \data_i[26][0] , \data_i[25][31] ,
         \data_i[25][30] , \data_i[25][29] , \data_i[25][28] ,
         \data_i[25][27] , \data_i[25][26] , \data_i[25][25] ,
         \data_i[25][24] , \data_i[25][23] , \data_i[25][22] ,
         \data_i[25][21] , \data_i[25][20] , \data_i[25][19] ,
         \data_i[25][18] , \data_i[25][17] , \data_i[25][16] ,
         \data_i[25][15] , \data_i[25][14] , \data_i[25][13] ,
         \data_i[25][12] , \data_i[25][11] , \data_i[25][10] , \data_i[25][9] ,
         \data_i[25][8] , \data_i[25][7] , \data_i[25][6] , \data_i[25][5] ,
         \data_i[25][4] , \data_i[25][3] , \data_i[25][2] , \data_i[25][1] ,
         \data_i[25][0] , \data_i[24][31] , \data_i[24][30] , \data_i[24][29] ,
         \data_i[24][28] , \data_i[24][27] , \data_i[24][26] ,
         \data_i[24][25] , \data_i[24][24] , \data_i[24][23] ,
         \data_i[24][22] , \data_i[24][21] , \data_i[24][20] ,
         \data_i[24][19] , \data_i[24][18] , \data_i[24][17] ,
         \data_i[24][16] , \data_i[24][15] , \data_i[24][14] ,
         \data_i[24][13] , \data_i[24][12] , \data_i[24][11] ,
         \data_i[24][10] , \data_i[24][9] , \data_i[24][8] , \data_i[24][7] ,
         \data_i[24][6] , \data_i[24][5] , \data_i[24][4] , \data_i[24][3] ,
         \data_i[24][2] , \data_i[24][1] , \data_i[24][0] , \data_i[23][31] ,
         \data_i[23][30] , \data_i[23][29] , \data_i[23][28] ,
         \data_i[23][27] , \data_i[23][26] , \data_i[23][25] ,
         \data_i[23][24] , \data_i[23][23] , \data_i[23][22] ,
         \data_i[23][21] , \data_i[23][20] , \data_i[23][19] ,
         \data_i[23][18] , \data_i[23][17] , \data_i[23][16] ,
         \data_i[23][15] , \data_i[23][14] , \data_i[23][13] ,
         \data_i[23][12] , \data_i[23][11] , \data_i[23][10] , \data_i[23][9] ,
         \data_i[23][8] , \data_i[23][7] , \data_i[23][6] , \data_i[23][5] ,
         \data_i[23][4] , \data_i[23][3] , \data_i[23][2] , \data_i[23][1] ,
         \data_i[23][0] , \data_i[22][31] , \data_i[22][30] , \data_i[22][29] ,
         \data_i[22][28] , \data_i[22][27] , \data_i[22][26] ,
         \data_i[22][25] , \data_i[22][24] , \data_i[22][23] ,
         \data_i[22][22] , \data_i[22][21] , \data_i[22][20] ,
         \data_i[22][19] , \data_i[22][18] , \data_i[22][17] ,
         \data_i[22][16] , \data_i[22][15] , \data_i[22][14] ,
         \data_i[22][13] , \data_i[22][12] , \data_i[22][11] ,
         \data_i[22][10] , \data_i[22][9] , \data_i[22][8] , \data_i[22][7] ,
         \data_i[22][6] , \data_i[22][5] , \data_i[22][4] , \data_i[22][3] ,
         \data_i[22][2] , \data_i[22][1] , \data_i[22][0] , \data_i[21][31] ,
         \data_i[21][30] , \data_i[21][29] , \data_i[21][28] ,
         \data_i[21][27] , \data_i[21][26] , \data_i[21][25] ,
         \data_i[21][24] , \data_i[21][23] , \data_i[21][22] ,
         \data_i[21][21] , \data_i[21][20] , \data_i[21][19] ,
         \data_i[21][18] , \data_i[21][17] , \data_i[21][16] ,
         \data_i[21][15] , \data_i[21][14] , \data_i[21][13] ,
         \data_i[21][12] , \data_i[21][11] , \data_i[21][10] , \data_i[21][9] ,
         \data_i[21][8] , \data_i[21][7] , \data_i[21][6] , \data_i[21][5] ,
         \data_i[21][4] , \data_i[21][3] , \data_i[21][2] , \data_i[21][1] ,
         \data_i[21][0] , \data_i[20][31] , \data_i[20][30] , \data_i[20][29] ,
         \data_i[20][28] , \data_i[20][27] , \data_i[20][26] ,
         \data_i[20][25] , \data_i[20][24] , \data_i[20][23] ,
         \data_i[20][22] , \data_i[20][21] , \data_i[20][20] ,
         \data_i[20][19] , \data_i[20][18] , \data_i[20][17] ,
         \data_i[20][16] , \data_i[20][15] , \data_i[20][14] ,
         \data_i[20][13] , \data_i[20][12] , \data_i[20][11] ,
         \data_i[20][10] , \data_i[20][9] , \data_i[20][8] , \data_i[20][7] ,
         \data_i[20][6] , \data_i[20][5] , \data_i[20][4] , \data_i[20][3] ,
         \data_i[20][2] , \data_i[20][1] , \data_i[20][0] , \data_i[19][31] ,
         \data_i[19][30] , \data_i[19][29] , \data_i[19][28] ,
         \data_i[19][27] , \data_i[19][26] , \data_i[19][25] ,
         \data_i[19][24] , \data_i[19][23] , \data_i[19][22] ,
         \data_i[19][21] , \data_i[19][20] , \data_i[19][19] ,
         \data_i[19][18] , \data_i[19][17] , \data_i[19][16] ,
         \data_i[19][15] , \data_i[19][14] , \data_i[19][13] ,
         \data_i[19][12] , \data_i[19][11] , \data_i[19][10] , \data_i[19][9] ,
         \data_i[19][8] , \data_i[19][7] , \data_i[19][6] , \data_i[19][5] ,
         \data_i[19][4] , \data_i[19][3] , \data_i[19][2] , \data_i[19][1] ,
         \data_i[19][0] , \data_i[18][31] , \data_i[18][30] , \data_i[18][29] ,
         \data_i[18][28] , \data_i[18][27] , \data_i[18][26] ,
         \data_i[18][25] , \data_i[18][24] , \data_i[18][23] ,
         \data_i[18][22] , \data_i[18][21] , \data_i[18][20] ,
         \data_i[18][19] , \data_i[18][18] , \data_i[18][17] ,
         \data_i[18][16] , \data_i[18][15] , \data_i[18][14] ,
         \data_i[18][13] , \data_i[18][12] , \data_i[18][11] ,
         \data_i[18][10] , \data_i[18][9] , \data_i[18][8] , \data_i[18][7] ,
         \data_i[18][6] , \data_i[18][5] , \data_i[18][4] , \data_i[18][3] ,
         \data_i[18][2] , \data_i[18][1] , \data_i[18][0] , \data_i[17][31] ,
         \data_i[17][30] , \data_i[17][29] , \data_i[17][28] ,
         \data_i[17][27] , \data_i[17][26] , \data_i[17][25] ,
         \data_i[17][24] , \data_i[17][23] , \data_i[17][22] ,
         \data_i[17][21] , \data_i[17][20] , \data_i[17][19] ,
         \data_i[17][18] , \data_i[17][17] , \data_i[17][16] ,
         \data_i[17][15] , \data_i[17][14] , \data_i[17][13] ,
         \data_i[17][12] , \data_i[17][11] , \data_i[17][10] , \data_i[17][9] ,
         \data_i[17][8] , \data_i[17][7] , \data_i[17][6] , \data_i[17][5] ,
         \data_i[17][4] , \data_i[17][3] , \data_i[17][2] , \data_i[17][1] ,
         \data_i[17][0] , \data_i[16][31] , \data_i[16][30] , \data_i[16][29] ,
         \data_i[16][28] , \data_i[16][27] , \data_i[16][26] ,
         \data_i[16][25] , \data_i[16][24] , \data_i[16][23] ,
         \data_i[16][22] , \data_i[16][21] , \data_i[16][20] ,
         \data_i[16][19] , \data_i[16][18] , \data_i[16][17] ,
         \data_i[16][16] , \data_i[16][15] , \data_i[16][14] ,
         \data_i[16][13] , \data_i[16][12] , \data_i[16][11] ,
         \data_i[16][10] , \data_i[16][9] , \data_i[16][8] , \data_i[16][7] ,
         \data_i[16][6] , \data_i[16][5] , \data_i[16][4] , \data_i[16][3] ,
         \data_i[16][2] , \data_i[16][1] , \data_i[16][0] , \data_i[15][31] ,
         \data_i[15][30] , \data_i[15][29] , \data_i[15][28] ,
         \data_i[15][27] , \data_i[15][26] , \data_i[15][25] ,
         \data_i[15][24] , \data_i[15][23] , \data_i[15][22] ,
         \data_i[15][21] , \data_i[15][20] , \data_i[15][19] ,
         \data_i[15][18] , \data_i[15][17] , \data_i[15][16] ,
         \data_i[15][15] , \data_i[15][14] , \data_i[15][13] ,
         \data_i[15][12] , \data_i[15][11] , \data_i[15][10] , \data_i[15][9] ,
         \data_i[15][8] , \data_i[15][7] , \data_i[15][6] , \data_i[15][5] ,
         \data_i[15][4] , \data_i[15][3] , \data_i[15][2] , \data_i[15][1] ,
         \data_i[15][0] , \data_i[14][31] , \data_i[14][30] , \data_i[14][29] ,
         \data_i[14][28] , \data_i[14][27] , \data_i[14][26] ,
         \data_i[14][25] , \data_i[14][24] , \data_i[14][23] ,
         \data_i[14][22] , \data_i[14][21] , \data_i[14][20] ,
         \data_i[14][19] , \data_i[14][18] , \data_i[14][17] ,
         \data_i[14][16] , \data_i[14][15] , \data_i[14][14] ,
         \data_i[14][13] , \data_i[14][12] , \data_i[14][11] ,
         \data_i[14][10] , \data_i[14][9] , \data_i[14][8] , \data_i[14][7] ,
         \data_i[14][6] , \data_i[14][5] , \data_i[14][4] , \data_i[14][3] ,
         \data_i[14][2] , \data_i[14][1] , \data_i[14][0] , \data_i[13][31] ,
         \data_i[13][30] , \data_i[13][29] , \data_i[13][28] ,
         \data_i[13][27] , \data_i[13][26] , \data_i[13][25] ,
         \data_i[13][24] , \data_i[13][23] , \data_i[13][22] ,
         \data_i[13][21] , \data_i[13][20] , \data_i[13][19] ,
         \data_i[13][18] , \data_i[13][17] , \data_i[13][16] ,
         \data_i[13][15] , \data_i[13][14] , \data_i[13][13] ,
         \data_i[13][12] , \data_i[13][11] , \data_i[13][10] , \data_i[13][9] ,
         \data_i[13][8] , \data_i[13][7] , \data_i[13][6] , \data_i[13][5] ,
         \data_i[13][4] , \data_i[13][3] , \data_i[13][2] , \data_i[13][1] ,
         \data_i[13][0] , \data_i[12][31] , \data_i[12][30] , \data_i[12][29] ,
         \data_i[12][28] , \data_i[12][27] , \data_i[12][26] ,
         \data_i[12][25] , \data_i[12][24] , \data_i[12][23] ,
         \data_i[12][22] , \data_i[12][21] , \data_i[12][20] ,
         \data_i[12][19] , \data_i[12][18] , \data_i[12][17] ,
         \data_i[12][16] , \data_i[12][15] , \data_i[12][14] ,
         \data_i[12][13] , \data_i[12][12] , \data_i[12][11] ,
         \data_i[12][10] , \data_i[12][9] , \data_i[12][8] , \data_i[12][7] ,
         \data_i[12][6] , \data_i[12][5] , \data_i[12][4] , \data_i[12][3] ,
         \data_i[12][2] , \data_i[12][1] , \data_i[12][0] , \data_i[11][31] ,
         \data_i[11][30] , \data_i[11][29] , \data_i[11][28] ,
         \data_i[11][27] , \data_i[11][26] , \data_i[11][25] ,
         \data_i[11][24] , \data_i[11][23] , \data_i[11][22] ,
         \data_i[11][21] , \data_i[11][20] , \data_i[11][19] ,
         \data_i[11][18] , \data_i[11][17] , \data_i[11][16] ,
         \data_i[11][15] , \data_i[11][14] , \data_i[11][13] ,
         \data_i[11][12] , \data_i[11][11] , \data_i[11][10] , \data_i[11][9] ,
         \data_i[11][8] , \data_i[11][7] , \data_i[11][6] , \data_i[11][5] ,
         \data_i[11][4] , \data_i[11][3] , \data_i[11][2] , \data_i[11][1] ,
         \data_i[11][0] , \data_i[10][31] , \data_i[10][30] , \data_i[10][29] ,
         \data_i[10][28] , \data_i[10][27] , \data_i[10][26] ,
         \data_i[10][25] , \data_i[10][24] , \data_i[10][23] ,
         \data_i[10][22] , \data_i[10][21] , \data_i[10][20] ,
         \data_i[10][19] , \data_i[10][18] , \data_i[10][17] ,
         \data_i[10][16] , \data_i[10][15] , \data_i[10][14] ,
         \data_i[10][13] , \data_i[10][12] , \data_i[10][11] ,
         \data_i[10][10] , \data_i[10][9] , \data_i[10][8] , \data_i[10][7] ,
         \data_i[10][6] , \data_i[10][5] , \data_i[10][4] , \data_i[10][3] ,
         \data_i[10][2] , \data_i[10][1] , \data_i[10][0] , \data_i[9][31] ,
         \data_i[9][30] , \data_i[9][29] , \data_i[9][28] , \data_i[9][27] ,
         \data_i[9][26] , \data_i[9][25] , \data_i[9][24] , \data_i[9][23] ,
         \data_i[9][22] , \data_i[9][21] , \data_i[9][20] , \data_i[9][19] ,
         \data_i[9][18] , \data_i[9][17] , \data_i[9][16] , \data_i[9][15] ,
         \data_i[9][14] , \data_i[9][13] , \data_i[9][12] , \data_i[9][11] ,
         \data_i[9][10] , \data_i[9][9] , \data_i[9][8] , \data_i[9][7] ,
         \data_i[9][6] , \data_i[9][5] , \data_i[9][4] , \data_i[9][3] ,
         \data_i[9][2] , \data_i[9][1] , \data_i[9][0] , \data_i[8][31] ,
         \data_i[8][30] , \data_i[8][29] , \data_i[8][28] , \data_i[8][27] ,
         \data_i[8][26] , \data_i[8][25] , \data_i[8][24] , \data_i[8][23] ,
         \data_i[8][22] , \data_i[8][21] , \data_i[8][20] , \data_i[8][19] ,
         \data_i[8][18] , \data_i[8][17] , \data_i[8][16] , \data_i[8][15] ,
         \data_i[8][14] , \data_i[8][13] , \data_i[8][12] , \data_i[8][11] ,
         \data_i[8][10] , \data_i[8][9] , \data_i[8][8] , \data_i[8][7] ,
         \data_i[8][6] , \data_i[8][5] , \data_i[8][4] , \data_i[8][3] ,
         \data_i[8][2] , \data_i[8][1] , \data_i[8][0] , \data_i[7][31] ,
         \data_i[7][30] , \data_i[7][29] , \data_i[7][28] , \data_i[7][27] ,
         \data_i[7][26] , \data_i[7][25] , \data_i[7][24] , \data_i[7][23] ,
         \data_i[7][22] , \data_i[7][21] , \data_i[7][20] , \data_i[7][19] ,
         \data_i[7][18] , \data_i[7][17] , \data_i[7][16] , \data_i[7][15] ,
         \data_i[7][14] , \data_i[7][13] , \data_i[7][12] , \data_i[7][11] ,
         \data_i[7][10] , \data_i[7][9] , \data_i[7][8] , \data_i[7][7] ,
         \data_i[7][6] , \data_i[7][5] , \data_i[7][4] , \data_i[7][3] ,
         \data_i[7][2] , \data_i[7][1] , \data_i[7][0] , \data_i[6][31] ,
         \data_i[6][30] , \data_i[6][29] , \data_i[6][28] , \data_i[6][27] ,
         \data_i[6][26] , \data_i[6][25] , \data_i[6][24] , \data_i[6][23] ,
         \data_i[6][22] , \data_i[6][21] , \data_i[6][20] , \data_i[6][19] ,
         \data_i[6][18] , \data_i[6][17] , \data_i[6][16] , \data_i[6][15] ,
         \data_i[6][14] , \data_i[6][13] , \data_i[6][12] , \data_i[6][11] ,
         \data_i[6][10] , \data_i[6][9] , \data_i[6][8] , \data_i[6][7] ,
         \data_i[6][6] , \data_i[6][5] , \data_i[6][4] , \data_i[6][3] ,
         \data_i[6][2] , \data_i[6][1] , \data_i[6][0] , \data_i[5][31] ,
         \data_i[5][30] , \data_i[5][29] , \data_i[5][28] , \data_i[5][27] ,
         \data_i[5][26] , \data_i[5][25] , \data_i[5][24] , \data_i[5][23] ,
         \data_i[5][22] , \data_i[5][21] , \data_i[5][20] , \data_i[5][19] ,
         \data_i[5][18] , \data_i[5][17] , \data_i[5][16] , \data_i[5][15] ,
         \data_i[5][14] , \data_i[5][13] , \data_i[5][12] , \data_i[5][11] ,
         \data_i[5][10] , \data_i[5][9] , \data_i[5][8] , \data_i[5][7] ,
         \data_i[5][6] , \data_i[5][5] , \data_i[5][4] , \data_i[5][3] ,
         \data_i[5][2] , \data_i[5][1] , \data_i[5][0] , \data_i[4][31] ,
         \data_i[4][30] , \data_i[4][29] , \data_i[4][28] , \data_i[4][27] ,
         \data_i[4][26] , \data_i[4][25] , \data_i[4][24] , \data_i[4][23] ,
         \data_i[4][22] , \data_i[4][21] , \data_i[4][20] , \data_i[4][19] ,
         \data_i[4][18] , \data_i[4][17] , \data_i[4][16] , \data_i[4][15] ,
         \data_i[4][14] , \data_i[4][13] , \data_i[4][12] , \data_i[4][11] ,
         \data_i[4][10] , \data_i[4][9] , \data_i[4][8] , \data_i[4][7] ,
         \data_i[4][6] , \data_i[4][5] , \data_i[4][4] , \data_i[4][3] ,
         \data_i[4][2] , \data_i[4][1] , \data_i[4][0] , \data_i[3][31] ,
         \data_i[3][30] , \data_i[3][29] , \data_i[3][28] , \data_i[3][27] ,
         \data_i[3][26] , \data_i[3][25] , \data_i[3][24] , \data_i[3][23] ,
         \data_i[3][22] , \data_i[3][21] , \data_i[3][20] , \data_i[3][19] ,
         \data_i[3][18] , \data_i[3][17] , \data_i[3][16] , \data_i[3][15] ,
         \data_i[3][14] , \data_i[3][13] , \data_i[3][12] , \data_i[3][11] ,
         \data_i[3][10] , \data_i[3][9] , \data_i[3][8] , \data_i[3][7] ,
         \data_i[3][6] , \data_i[3][5] , \data_i[3][4] , \data_i[3][3] ,
         \data_i[3][2] , \data_i[3][1] , \data_i[3][0] , \data_i[2][31] ,
         \data_i[2][30] , \data_i[2][29] , \data_i[2][28] , \data_i[2][27] ,
         \data_i[2][26] , \data_i[2][25] , \data_i[2][24] , \data_i[2][23] ,
         \data_i[2][22] , \data_i[2][21] , \data_i[2][20] , \data_i[2][19] ,
         \data_i[2][18] , \data_i[2][17] , \data_i[2][16] , \data_i[2][15] ,
         \data_i[2][14] , \data_i[2][13] , \data_i[2][12] , \data_i[2][11] ,
         \data_i[2][10] , \data_i[2][9] , \data_i[2][8] , \data_i[2][7] ,
         \data_i[2][6] , \data_i[2][5] , \data_i[2][4] , \data_i[2][3] ,
         \data_i[2][2] , \data_i[2][1] , \data_i[2][0] , \data_i[1][31] ,
         \data_i[1][30] , \data_i[1][29] , \data_i[1][28] , \data_i[1][27] ,
         \data_i[1][26] , \data_i[1][25] , \data_i[1][24] , \data_i[1][23] ,
         \data_i[1][22] , \data_i[1][21] , \data_i[1][20] , \data_i[1][19] ,
         \data_i[1][18] , \data_i[1][17] , \data_i[1][16] , \data_i[1][15] ,
         \data_i[1][14] , \data_i[1][13] , \data_i[1][12] , \data_i[1][11] ,
         \data_i[1][10] , \data_i[1][9] , \data_i[1][8] , \data_i[1][7] ,
         \data_i[1][6] , \data_i[1][5] , \data_i[1][4] , \data_i[1][3] ,
         \data_i[1][2] , \data_i[1][1] , \data_i[1][0] , \data_i[0][31] ,
         \data_i[0][30] , \data_i[0][29] , \data_i[0][28] , \data_i[0][27] ,
         \data_i[0][26] , \data_i[0][25] , \data_i[0][24] , \data_i[0][23] ,
         \data_i[0][22] , \data_i[0][21] , \data_i[0][20] , \data_i[0][19] ,
         \data_i[0][18] , \data_i[0][17] , \data_i[0][16] , \data_i[0][15] ,
         \data_i[0][14] , \data_i[0][13] , \data_i[0][12] , \data_i[0][11] ,
         \data_i[0][10] , \data_i[0][9] , \data_i[0][8] , \data_i[0][7] ,
         \data_i[0][6] , \data_i[0][5] , \data_i[0][4] , \data_i[0][3] ,
         \data_i[0][2] , \data_i[0][1] , \data_i[0][0] ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698;

  INVD1 U1 ( .I(select_i[4]), .ZN(n645) );
  INVD1 U2 ( .I(select_i[2]), .ZN(n641) );
  NR2D1 U3 ( .A1(select_i[2]), .A2(n650), .ZN(n652) );
  INVD1 U4 ( .I(select_i[3]), .ZN(n651) );
  INVD1 U5 ( .I(select_i[1]), .ZN(n650) );
  INVD1 U6 ( .I(select_i[0]), .ZN(n643) );
  NR2D1 U7 ( .A1(select_i[3]), .A2(n641), .ZN(n642) );
  ND2D1 U8 ( .A1(select_i[3]), .A2(n645), .ZN(n647) );
  ND2D1 U9 ( .A1(n652), .A2(n645), .ZN(n646) );
  OR2XD1 U10 ( .A1(n648), .A2(select_i[2]), .Z(n644) );
  ND2D1 U11 ( .A1(n645), .A2(n650), .ZN(n648) );
  ND2D1 U12 ( .A1(select_i[1]), .A2(n645), .ZN(n649) );
  IND2D1 U13 ( .A1(n660), .B1(select_i[2]), .ZN(n664) );
  ND3D1 U14 ( .A1(select_i[2]), .A2(select_i[3]), .A3(select_i[0]), .ZN(n666)
         );
  ND2D1 U15 ( .A1(select_i[3]), .A2(n643), .ZN(n660) );
  ND2D1 U16 ( .A1(select_i[4]), .A2(select_i[3]), .ZN(n661) );
  OR2XD1 U17 ( .A1(n663), .A2(select_i[2]), .Z(n657) );
  ND3D1 U18 ( .A1(select_i[0]), .A2(n641), .A3(n650), .ZN(n658) );
  ND2D1 U19 ( .A1(n651), .A2(n643), .ZN(n653) );
  ND2D1 U20 ( .A1(select_i[0]), .A2(n652), .ZN(n662) );
  ND2D1 U21 ( .A1(select_i[4]), .A2(n651), .ZN(n654) );
  ND2D1 U22 ( .A1(select_i[4]), .A2(select_i[1]), .ZN(n665) );
  ND2D1 U23 ( .A1(select_i[0]), .A2(n642), .ZN(n656) );
  ND2D1 U24 ( .A1(n650), .A2(select_i[4]), .ZN(n663) );
  ND2D1 U25 ( .A1(n642), .A2(n643), .ZN(n655) );
  NR2D1 U26 ( .A1(n649), .A2(n664), .ZN(n682) );
  NR2D1 U27 ( .A1(n649), .A2(n666), .ZN(n681) );
  NR2D1 U28 ( .A1(n648), .A2(n664), .ZN(n680) );
  NR2D1 U29 ( .A1(n648), .A2(n666), .ZN(n679) );
  NR2D1 U30 ( .A1(n644), .A2(n660), .ZN(n676) );
  NR2D1 U31 ( .A1(n658), .A2(n647), .ZN(n675) );
  NR2D1 U32 ( .A1(n662), .A2(n647), .ZN(n677) );
  NR2D1 U33 ( .A1(n646), .A2(n660), .ZN(n678) );
  NR3D1 U34 ( .A1(select_i[4]), .A2(select_i[3]), .A3(n662), .ZN(n669) );
  NR2D1 U35 ( .A1(n653), .A2(n646), .ZN(n670) );
  NR2D1 U36 ( .A1(n644), .A2(n653), .ZN(n668) );
  NR3D1 U37 ( .A1(select_i[4]), .A2(select_i[3]), .A3(n658), .ZN(n667) );
  NR2D1 U38 ( .A1(n648), .A2(n656), .ZN(n671) );
  NR2D1 U39 ( .A1(n648), .A2(n655), .ZN(n672) );
  NR2D1 U40 ( .A1(n656), .A2(n649), .ZN(n673) );
  NR2D1 U41 ( .A1(n655), .A2(n649), .ZN(n674) );
  NR2D1 U42 ( .A1(n664), .A2(n665), .ZN(n698) );
  NR2D1 U43 ( .A1(n666), .A2(n665), .ZN(n697) );
  NR2D1 U44 ( .A1(n664), .A2(n663), .ZN(n696) );
  NR2D1 U45 ( .A1(n666), .A2(n663), .ZN(n695) );
  NR2D1 U46 ( .A1(n660), .A2(n657), .ZN(n692) );
  NR2D1 U47 ( .A1(n658), .A2(n661), .ZN(n691) );
  NR2D1 U48 ( .A1(n660), .A2(n659), .ZN(n694) );
  NR2D1 U49 ( .A1(n662), .A2(n661), .ZN(n693) );
  NR2D1 U50 ( .A1(n653), .A2(n657), .ZN(n684) );
  NR2D1 U51 ( .A1(n658), .A2(n654), .ZN(n683) );
  NR2D1 U52 ( .A1(n653), .A2(n659), .ZN(n686) );
  NR2D1 U53 ( .A1(n662), .A2(n654), .ZN(n685) );
  NR2D1 U54 ( .A1(n656), .A2(n665), .ZN(n689) );
  NR2D1 U55 ( .A1(n655), .A2(n665), .ZN(n690) );
  NR2D1 U56 ( .A1(n656), .A2(n663), .ZN(n687) );
  NR2D1 U57 ( .A1(n655), .A2(n663), .ZN(n688) );
  AOI22D0 U58 ( .A1(\data_i[17][0] ), .A2(n683), .B1(\data_i[16][0] ), .B2(
        n684), .ZN(n1) );
  AOI22D0 U59 ( .A1(\data_i[19][0] ), .A2(n685), .B1(\data_i[18][0] ), .B2(
        n686), .ZN(n2) );
  AOI22D0 U60 ( .A1(\data_i[21][0] ), .A2(n687), .B1(\data_i[20][0] ), .B2(
        n688), .ZN(n3) );
  AOI22D0 U61 ( .A1(\data_i[23][0] ), .A2(n689), .B1(\data_i[22][0] ), .B2(
        n690), .ZN(n4) );
  ND4D0 U62 ( .A1(n1), .A2(n2), .A3(n3), .A4(n4), .ZN(n5) );
  AOI22D0 U63 ( .A1(\data_i[25][0] ), .A2(n691), .B1(\data_i[24][0] ), .B2(
        n692), .ZN(n6) );
  AOI22D0 U64 ( .A1(\data_i[27][0] ), .A2(n693), .B1(\data_i[26][0] ), .B2(
        n694), .ZN(n7) );
  AOI22D0 U65 ( .A1(\data_i[29][0] ), .A2(n695), .B1(\data_i[28][0] ), .B2(
        n696), .ZN(n8) );
  AOI22D0 U66 ( .A1(\data_i[31][0] ), .A2(n697), .B1(\data_i[30][0] ), .B2(
        n698), .ZN(n9) );
  ND4D0 U67 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .ZN(n10) );
  AOI22D0 U68 ( .A1(\data_i[1][0] ), .A2(n667), .B1(\data_i[0][0] ), .B2(n668), 
        .ZN(n11) );
  AOI22D0 U69 ( .A1(\data_i[3][0] ), .A2(n669), .B1(\data_i[2][0] ), .B2(n670), 
        .ZN(n12) );
  AOI22D0 U70 ( .A1(\data_i[5][0] ), .A2(n671), .B1(\data_i[4][0] ), .B2(n672), 
        .ZN(n13) );
  AOI22D0 U71 ( .A1(\data_i[7][0] ), .A2(n673), .B1(\data_i[6][0] ), .B2(n674), 
        .ZN(n14) );
  ND4D0 U72 ( .A1(n11), .A2(n12), .A3(n13), .A4(n14), .ZN(n15) );
  AOI22D0 U73 ( .A1(\data_i[9][0] ), .A2(n675), .B1(\data_i[8][0] ), .B2(n676), 
        .ZN(n16) );
  AOI22D0 U74 ( .A1(\data_i[11][0] ), .A2(n677), .B1(\data_i[10][0] ), .B2(
        n678), .ZN(n17) );
  AOI22D0 U75 ( .A1(\data_i[13][0] ), .A2(n679), .B1(\data_i[12][0] ), .B2(
        n680), .ZN(n18) );
  AOI22D0 U76 ( .A1(\data_i[15][0] ), .A2(n681), .B1(\data_i[14][0] ), .B2(
        n682), .ZN(n19) );
  ND4D0 U77 ( .A1(n16), .A2(n17), .A3(n18), .A4(n19), .ZN(n20) );
  OR4D0 U78 ( .A1(n5), .A2(n10), .A3(n15), .A4(n20), .Z(data_o[0]) );
  AOI22D0 U79 ( .A1(\data_i[17][1] ), .A2(n683), .B1(\data_i[16][1] ), .B2(
        n684), .ZN(n21) );
  AOI22D0 U80 ( .A1(\data_i[19][1] ), .A2(n685), .B1(\data_i[18][1] ), .B2(
        n686), .ZN(n22) );
  AOI22D0 U81 ( .A1(\data_i[21][1] ), .A2(n687), .B1(\data_i[20][1] ), .B2(
        n688), .ZN(n23) );
  AOI22D0 U82 ( .A1(\data_i[23][1] ), .A2(n689), .B1(\data_i[22][1] ), .B2(
        n690), .ZN(n24) );
  ND4D0 U83 ( .A1(n21), .A2(n22), .A3(n23), .A4(n24), .ZN(n25) );
  AOI22D0 U84 ( .A1(\data_i[25][1] ), .A2(n691), .B1(\data_i[24][1] ), .B2(
        n692), .ZN(n26) );
  AOI22D0 U85 ( .A1(\data_i[27][1] ), .A2(n693), .B1(\data_i[26][1] ), .B2(
        n694), .ZN(n27) );
  AOI22D0 U86 ( .A1(\data_i[29][1] ), .A2(n695), .B1(\data_i[28][1] ), .B2(
        n696), .ZN(n28) );
  AOI22D0 U87 ( .A1(\data_i[31][1] ), .A2(n697), .B1(\data_i[30][1] ), .B2(
        n698), .ZN(n29) );
  ND4D0 U88 ( .A1(n26), .A2(n27), .A3(n28), .A4(n29), .ZN(n30) );
  AOI22D0 U89 ( .A1(\data_i[1][1] ), .A2(n667), .B1(\data_i[0][1] ), .B2(n668), 
        .ZN(n31) );
  AOI22D0 U90 ( .A1(\data_i[3][1] ), .A2(n669), .B1(\data_i[2][1] ), .B2(n670), 
        .ZN(n32) );
  AOI22D0 U91 ( .A1(\data_i[5][1] ), .A2(n671), .B1(\data_i[4][1] ), .B2(n672), 
        .ZN(n33) );
  AOI22D0 U92 ( .A1(\data_i[7][1] ), .A2(n673), .B1(\data_i[6][1] ), .B2(n674), 
        .ZN(n34) );
  ND4D0 U93 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(n35) );
  AOI22D0 U94 ( .A1(\data_i[9][1] ), .A2(n675), .B1(\data_i[8][1] ), .B2(n676), 
        .ZN(n36) );
  AOI22D0 U95 ( .A1(\data_i[11][1] ), .A2(n677), .B1(\data_i[10][1] ), .B2(
        n678), .ZN(n37) );
  AOI22D0 U96 ( .A1(\data_i[13][1] ), .A2(n679), .B1(\data_i[12][1] ), .B2(
        n680), .ZN(n38) );
  AOI22D0 U97 ( .A1(\data_i[15][1] ), .A2(n681), .B1(\data_i[14][1] ), .B2(
        n682), .ZN(n39) );
  ND4D0 U98 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .ZN(n40) );
  OR4D0 U99 ( .A1(n25), .A2(n30), .A3(n35), .A4(n40), .Z(data_o[1]) );
  AOI22D0 U100 ( .A1(\data_i[17][2] ), .A2(n683), .B1(\data_i[16][2] ), .B2(
        n684), .ZN(n41) );
  AOI22D0 U101 ( .A1(\data_i[19][2] ), .A2(n685), .B1(\data_i[18][2] ), .B2(
        n686), .ZN(n42) );
  AOI22D0 U102 ( .A1(\data_i[21][2] ), .A2(n687), .B1(\data_i[20][2] ), .B2(
        n688), .ZN(n43) );
  AOI22D0 U103 ( .A1(\data_i[23][2] ), .A2(n689), .B1(\data_i[22][2] ), .B2(
        n690), .ZN(n44) );
  ND4D0 U104 ( .A1(n41), .A2(n42), .A3(n43), .A4(n44), .ZN(n45) );
  AOI22D0 U105 ( .A1(\data_i[25][2] ), .A2(n691), .B1(\data_i[24][2] ), .B2(
        n692), .ZN(n46) );
  AOI22D0 U106 ( .A1(\data_i[27][2] ), .A2(n693), .B1(\data_i[26][2] ), .B2(
        n694), .ZN(n47) );
  AOI22D0 U107 ( .A1(\data_i[29][2] ), .A2(n695), .B1(\data_i[28][2] ), .B2(
        n696), .ZN(n48) );
  AOI22D0 U108 ( .A1(\data_i[31][2] ), .A2(n697), .B1(\data_i[30][2] ), .B2(
        n698), .ZN(n49) );
  ND4D0 U109 ( .A1(n46), .A2(n47), .A3(n48), .A4(n49), .ZN(n50) );
  AOI22D0 U110 ( .A1(\data_i[1][2] ), .A2(n667), .B1(\data_i[0][2] ), .B2(n668), .ZN(n51) );
  AOI22D0 U111 ( .A1(\data_i[3][2] ), .A2(n669), .B1(\data_i[2][2] ), .B2(n670), .ZN(n52) );
  AOI22D0 U112 ( .A1(\data_i[5][2] ), .A2(n671), .B1(\data_i[4][2] ), .B2(n672), .ZN(n53) );
  AOI22D0 U113 ( .A1(\data_i[7][2] ), .A2(n673), .B1(\data_i[6][2] ), .B2(n674), .ZN(n54) );
  ND4D0 U114 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(n55) );
  AOI22D0 U115 ( .A1(\data_i[9][2] ), .A2(n675), .B1(\data_i[8][2] ), .B2(n676), .ZN(n56) );
  AOI22D0 U116 ( .A1(\data_i[11][2] ), .A2(n677), .B1(\data_i[10][2] ), .B2(
        n678), .ZN(n57) );
  AOI22D0 U117 ( .A1(\data_i[13][2] ), .A2(n679), .B1(\data_i[12][2] ), .B2(
        n680), .ZN(n58) );
  AOI22D0 U118 ( .A1(\data_i[15][2] ), .A2(n681), .B1(\data_i[14][2] ), .B2(
        n682), .ZN(n59) );
  ND4D0 U119 ( .A1(n56), .A2(n57), .A3(n58), .A4(n59), .ZN(n60) );
  OR4D0 U120 ( .A1(n45), .A2(n50), .A3(n55), .A4(n60), .Z(data_o[2]) );
  AOI22D0 U121 ( .A1(\data_i[17][3] ), .A2(n683), .B1(\data_i[16][3] ), .B2(
        n684), .ZN(n61) );
  AOI22D0 U122 ( .A1(\data_i[19][3] ), .A2(n685), .B1(\data_i[18][3] ), .B2(
        n686), .ZN(n62) );
  AOI22D0 U123 ( .A1(\data_i[21][3] ), .A2(n687), .B1(\data_i[20][3] ), .B2(
        n688), .ZN(n63) );
  AOI22D0 U124 ( .A1(\data_i[23][3] ), .A2(n689), .B1(\data_i[22][3] ), .B2(
        n690), .ZN(n64) );
  ND4D0 U125 ( .A1(n61), .A2(n62), .A3(n63), .A4(n64), .ZN(n65) );
  AOI22D0 U126 ( .A1(\data_i[25][3] ), .A2(n691), .B1(\data_i[24][3] ), .B2(
        n692), .ZN(n66) );
  AOI22D0 U127 ( .A1(\data_i[27][3] ), .A2(n693), .B1(\data_i[26][3] ), .B2(
        n694), .ZN(n67) );
  AOI22D0 U128 ( .A1(\data_i[29][3] ), .A2(n695), .B1(\data_i[28][3] ), .B2(
        n696), .ZN(n68) );
  AOI22D0 U129 ( .A1(\data_i[31][3] ), .A2(n697), .B1(\data_i[30][3] ), .B2(
        n698), .ZN(n69) );
  ND4D0 U130 ( .A1(n66), .A2(n67), .A3(n68), .A4(n69), .ZN(n70) );
  AOI22D0 U131 ( .A1(\data_i[1][3] ), .A2(n667), .B1(\data_i[0][3] ), .B2(n668), .ZN(n71) );
  AOI22D0 U132 ( .A1(\data_i[3][3] ), .A2(n669), .B1(\data_i[2][3] ), .B2(n670), .ZN(n72) );
  AOI22D0 U133 ( .A1(\data_i[5][3] ), .A2(n671), .B1(\data_i[4][3] ), .B2(n672), .ZN(n73) );
  AOI22D0 U134 ( .A1(\data_i[7][3] ), .A2(n673), .B1(\data_i[6][3] ), .B2(n674), .ZN(n74) );
  ND4D0 U135 ( .A1(n71), .A2(n72), .A3(n73), .A4(n74), .ZN(n75) );
  AOI22D0 U136 ( .A1(\data_i[9][3] ), .A2(n675), .B1(\data_i[8][3] ), .B2(n676), .ZN(n76) );
  AOI22D0 U137 ( .A1(\data_i[11][3] ), .A2(n677), .B1(\data_i[10][3] ), .B2(
        n678), .ZN(n77) );
  AOI22D0 U138 ( .A1(\data_i[13][3] ), .A2(n679), .B1(\data_i[12][3] ), .B2(
        n680), .ZN(n78) );
  AOI22D0 U139 ( .A1(\data_i[15][3] ), .A2(n681), .B1(\data_i[14][3] ), .B2(
        n682), .ZN(n79) );
  ND4D0 U140 ( .A1(n76), .A2(n77), .A3(n78), .A4(n79), .ZN(n80) );
  OR4D0 U141 ( .A1(n65), .A2(n70), .A3(n75), .A4(n80), .Z(data_o[3]) );
  AOI22D0 U142 ( .A1(\data_i[17][4] ), .A2(n683), .B1(\data_i[16][4] ), .B2(
        n684), .ZN(n81) );
  AOI22D0 U143 ( .A1(\data_i[19][4] ), .A2(n685), .B1(\data_i[18][4] ), .B2(
        n686), .ZN(n82) );
  AOI22D0 U144 ( .A1(\data_i[21][4] ), .A2(n687), .B1(\data_i[20][4] ), .B2(
        n688), .ZN(n83) );
  AOI22D0 U145 ( .A1(\data_i[23][4] ), .A2(n689), .B1(\data_i[22][4] ), .B2(
        n690), .ZN(n84) );
  ND4D0 U146 ( .A1(n81), .A2(n82), .A3(n83), .A4(n84), .ZN(n85) );
  AOI22D0 U147 ( .A1(\data_i[25][4] ), .A2(n691), .B1(\data_i[24][4] ), .B2(
        n692), .ZN(n86) );
  AOI22D0 U148 ( .A1(\data_i[27][4] ), .A2(n693), .B1(\data_i[26][4] ), .B2(
        n694), .ZN(n87) );
  AOI22D0 U149 ( .A1(\data_i[29][4] ), .A2(n695), .B1(\data_i[28][4] ), .B2(
        n696), .ZN(n88) );
  AOI22D0 U150 ( .A1(\data_i[31][4] ), .A2(n697), .B1(\data_i[30][4] ), .B2(
        n698), .ZN(n89) );
  ND4D0 U151 ( .A1(n86), .A2(n87), .A3(n88), .A4(n89), .ZN(n90) );
  AOI22D0 U152 ( .A1(\data_i[1][4] ), .A2(n667), .B1(\data_i[0][4] ), .B2(n668), .ZN(n91) );
  AOI22D0 U153 ( .A1(\data_i[3][4] ), .A2(n669), .B1(\data_i[2][4] ), .B2(n670), .ZN(n92) );
  AOI22D0 U154 ( .A1(\data_i[5][4] ), .A2(n671), .B1(\data_i[4][4] ), .B2(n672), .ZN(n93) );
  AOI22D0 U155 ( .A1(\data_i[7][4] ), .A2(n673), .B1(\data_i[6][4] ), .B2(n674), .ZN(n94) );
  ND4D0 U156 ( .A1(n91), .A2(n92), .A3(n93), .A4(n94), .ZN(n95) );
  AOI22D0 U157 ( .A1(\data_i[9][4] ), .A2(n675), .B1(\data_i[8][4] ), .B2(n676), .ZN(n96) );
  AOI22D0 U158 ( .A1(\data_i[11][4] ), .A2(n677), .B1(\data_i[10][4] ), .B2(
        n678), .ZN(n97) );
  AOI22D0 U159 ( .A1(\data_i[13][4] ), .A2(n679), .B1(\data_i[12][4] ), .B2(
        n680), .ZN(n98) );
  AOI22D0 U160 ( .A1(\data_i[15][4] ), .A2(n681), .B1(\data_i[14][4] ), .B2(
        n682), .ZN(n99) );
  ND4D0 U161 ( .A1(n96), .A2(n97), .A3(n98), .A4(n99), .ZN(n100) );
  OR4D0 U162 ( .A1(n85), .A2(n90), .A3(n95), .A4(n100), .Z(data_o[4]) );
  AOI22D0 U163 ( .A1(\data_i[17][5] ), .A2(n683), .B1(\data_i[16][5] ), .B2(
        n684), .ZN(n101) );
  AOI22D0 U164 ( .A1(\data_i[19][5] ), .A2(n685), .B1(\data_i[18][5] ), .B2(
        n686), .ZN(n102) );
  AOI22D0 U165 ( .A1(\data_i[21][5] ), .A2(n687), .B1(\data_i[20][5] ), .B2(
        n688), .ZN(n103) );
  AOI22D0 U166 ( .A1(\data_i[23][5] ), .A2(n689), .B1(\data_i[22][5] ), .B2(
        n690), .ZN(n104) );
  ND4D0 U167 ( .A1(n101), .A2(n102), .A3(n103), .A4(n104), .ZN(n105) );
  AOI22D0 U168 ( .A1(\data_i[25][5] ), .A2(n691), .B1(\data_i[24][5] ), .B2(
        n692), .ZN(n106) );
  AOI22D0 U169 ( .A1(\data_i[27][5] ), .A2(n693), .B1(\data_i[26][5] ), .B2(
        n694), .ZN(n107) );
  AOI22D0 U170 ( .A1(\data_i[29][5] ), .A2(n695), .B1(\data_i[28][5] ), .B2(
        n696), .ZN(n108) );
  AOI22D0 U171 ( .A1(\data_i[31][5] ), .A2(n697), .B1(\data_i[30][5] ), .B2(
        n698), .ZN(n109) );
  ND4D0 U172 ( .A1(n106), .A2(n107), .A3(n108), .A4(n109), .ZN(n110) );
  AOI22D0 U173 ( .A1(\data_i[1][5] ), .A2(n667), .B1(\data_i[0][5] ), .B2(n668), .ZN(n111) );
  AOI22D0 U174 ( .A1(\data_i[3][5] ), .A2(n669), .B1(\data_i[2][5] ), .B2(n670), .ZN(n112) );
  AOI22D0 U175 ( .A1(\data_i[5][5] ), .A2(n671), .B1(\data_i[4][5] ), .B2(n672), .ZN(n113) );
  AOI22D0 U176 ( .A1(\data_i[7][5] ), .A2(n673), .B1(\data_i[6][5] ), .B2(n674), .ZN(n114) );
  ND4D0 U177 ( .A1(n111), .A2(n112), .A3(n113), .A4(n114), .ZN(n115) );
  AOI22D0 U178 ( .A1(\data_i[9][5] ), .A2(n675), .B1(\data_i[8][5] ), .B2(n676), .ZN(n116) );
  AOI22D0 U179 ( .A1(\data_i[11][5] ), .A2(n677), .B1(\data_i[10][5] ), .B2(
        n678), .ZN(n117) );
  AOI22D0 U180 ( .A1(\data_i[13][5] ), .A2(n679), .B1(\data_i[12][5] ), .B2(
        n680), .ZN(n118) );
  AOI22D0 U181 ( .A1(\data_i[15][5] ), .A2(n681), .B1(\data_i[14][5] ), .B2(
        n682), .ZN(n119) );
  ND4D0 U182 ( .A1(n116), .A2(n117), .A3(n118), .A4(n119), .ZN(n120) );
  OR4D0 U183 ( .A1(n105), .A2(n110), .A3(n115), .A4(n120), .Z(data_o[5]) );
  AOI22D0 U184 ( .A1(\data_i[17][6] ), .A2(n683), .B1(\data_i[16][6] ), .B2(
        n684), .ZN(n121) );
  AOI22D0 U185 ( .A1(\data_i[19][6] ), .A2(n685), .B1(\data_i[18][6] ), .B2(
        n686), .ZN(n122) );
  AOI22D0 U186 ( .A1(\data_i[21][6] ), .A2(n687), .B1(\data_i[20][6] ), .B2(
        n688), .ZN(n123) );
  AOI22D0 U187 ( .A1(\data_i[23][6] ), .A2(n689), .B1(\data_i[22][6] ), .B2(
        n690), .ZN(n124) );
  ND4D0 U188 ( .A1(n121), .A2(n122), .A3(n123), .A4(n124), .ZN(n125) );
  AOI22D0 U189 ( .A1(\data_i[25][6] ), .A2(n691), .B1(\data_i[24][6] ), .B2(
        n692), .ZN(n126) );
  AOI22D0 U190 ( .A1(\data_i[27][6] ), .A2(n693), .B1(\data_i[26][6] ), .B2(
        n694), .ZN(n127) );
  AOI22D0 U191 ( .A1(\data_i[29][6] ), .A2(n695), .B1(\data_i[28][6] ), .B2(
        n696), .ZN(n128) );
  AOI22D0 U192 ( .A1(\data_i[31][6] ), .A2(n697), .B1(\data_i[30][6] ), .B2(
        n698), .ZN(n129) );
  ND4D0 U193 ( .A1(n126), .A2(n127), .A3(n128), .A4(n129), .ZN(n130) );
  AOI22D0 U194 ( .A1(\data_i[1][6] ), .A2(n667), .B1(\data_i[0][6] ), .B2(n668), .ZN(n131) );
  AOI22D0 U195 ( .A1(\data_i[3][6] ), .A2(n669), .B1(\data_i[2][6] ), .B2(n670), .ZN(n132) );
  AOI22D0 U196 ( .A1(\data_i[5][6] ), .A2(n671), .B1(\data_i[4][6] ), .B2(n672), .ZN(n133) );
  AOI22D0 U197 ( .A1(\data_i[7][6] ), .A2(n673), .B1(\data_i[6][6] ), .B2(n674), .ZN(n134) );
  ND4D0 U198 ( .A1(n131), .A2(n132), .A3(n133), .A4(n134), .ZN(n135) );
  AOI22D0 U199 ( .A1(\data_i[9][6] ), .A2(n675), .B1(\data_i[8][6] ), .B2(n676), .ZN(n136) );
  AOI22D0 U200 ( .A1(\data_i[11][6] ), .A2(n677), .B1(\data_i[10][6] ), .B2(
        n678), .ZN(n137) );
  AOI22D0 U201 ( .A1(\data_i[13][6] ), .A2(n679), .B1(\data_i[12][6] ), .B2(
        n680), .ZN(n138) );
  AOI22D0 U202 ( .A1(\data_i[15][6] ), .A2(n681), .B1(\data_i[14][6] ), .B2(
        n682), .ZN(n139) );
  ND4D0 U203 ( .A1(n136), .A2(n137), .A3(n138), .A4(n139), .ZN(n140) );
  OR4D0 U204 ( .A1(n125), .A2(n130), .A3(n135), .A4(n140), .Z(data_o[6]) );
  AOI22D0 U205 ( .A1(\data_i[17][7] ), .A2(n683), .B1(\data_i[16][7] ), .B2(
        n684), .ZN(n141) );
  AOI22D0 U206 ( .A1(\data_i[19][7] ), .A2(n685), .B1(\data_i[18][7] ), .B2(
        n686), .ZN(n142) );
  AOI22D0 U207 ( .A1(\data_i[21][7] ), .A2(n687), .B1(\data_i[20][7] ), .B2(
        n688), .ZN(n143) );
  AOI22D0 U208 ( .A1(\data_i[23][7] ), .A2(n689), .B1(\data_i[22][7] ), .B2(
        n690), .ZN(n144) );
  ND4D0 U209 ( .A1(n141), .A2(n142), .A3(n143), .A4(n144), .ZN(n145) );
  AOI22D0 U210 ( .A1(\data_i[25][7] ), .A2(n691), .B1(\data_i[24][7] ), .B2(
        n692), .ZN(n146) );
  AOI22D0 U211 ( .A1(\data_i[27][7] ), .A2(n693), .B1(\data_i[26][7] ), .B2(
        n694), .ZN(n147) );
  AOI22D0 U212 ( .A1(\data_i[29][7] ), .A2(n695), .B1(\data_i[28][7] ), .B2(
        n696), .ZN(n148) );
  AOI22D0 U213 ( .A1(\data_i[31][7] ), .A2(n697), .B1(\data_i[30][7] ), .B2(
        n698), .ZN(n149) );
  ND4D0 U214 ( .A1(n146), .A2(n147), .A3(n148), .A4(n149), .ZN(n150) );
  AOI22D0 U215 ( .A1(\data_i[1][7] ), .A2(n667), .B1(\data_i[0][7] ), .B2(n668), .ZN(n151) );
  AOI22D0 U216 ( .A1(\data_i[3][7] ), .A2(n669), .B1(\data_i[2][7] ), .B2(n670), .ZN(n152) );
  AOI22D0 U217 ( .A1(\data_i[5][7] ), .A2(n671), .B1(\data_i[4][7] ), .B2(n672), .ZN(n153) );
  AOI22D0 U218 ( .A1(\data_i[7][7] ), .A2(n673), .B1(\data_i[6][7] ), .B2(n674), .ZN(n154) );
  ND4D0 U219 ( .A1(n151), .A2(n152), .A3(n153), .A4(n154), .ZN(n155) );
  AOI22D0 U220 ( .A1(\data_i[9][7] ), .A2(n675), .B1(\data_i[8][7] ), .B2(n676), .ZN(n156) );
  AOI22D0 U221 ( .A1(\data_i[11][7] ), .A2(n677), .B1(\data_i[10][7] ), .B2(
        n678), .ZN(n157) );
  AOI22D0 U222 ( .A1(\data_i[13][7] ), .A2(n679), .B1(\data_i[12][7] ), .B2(
        n680), .ZN(n158) );
  AOI22D0 U223 ( .A1(\data_i[15][7] ), .A2(n681), .B1(\data_i[14][7] ), .B2(
        n682), .ZN(n159) );
  ND4D0 U224 ( .A1(n156), .A2(n157), .A3(n158), .A4(n159), .ZN(n160) );
  OR4D0 U225 ( .A1(n145), .A2(n150), .A3(n155), .A4(n160), .Z(data_o[7]) );
  AOI22D0 U226 ( .A1(\data_i[17][8] ), .A2(n683), .B1(\data_i[16][8] ), .B2(
        n684), .ZN(n161) );
  AOI22D0 U227 ( .A1(\data_i[19][8] ), .A2(n685), .B1(\data_i[18][8] ), .B2(
        n686), .ZN(n162) );
  AOI22D0 U228 ( .A1(\data_i[21][8] ), .A2(n687), .B1(\data_i[20][8] ), .B2(
        n688), .ZN(n163) );
  AOI22D0 U229 ( .A1(\data_i[23][8] ), .A2(n689), .B1(\data_i[22][8] ), .B2(
        n690), .ZN(n164) );
  ND4D0 U230 ( .A1(n161), .A2(n162), .A3(n163), .A4(n164), .ZN(n165) );
  AOI22D0 U231 ( .A1(\data_i[25][8] ), .A2(n691), .B1(\data_i[24][8] ), .B2(
        n692), .ZN(n166) );
  AOI22D0 U232 ( .A1(\data_i[27][8] ), .A2(n693), .B1(\data_i[26][8] ), .B2(
        n694), .ZN(n167) );
  AOI22D0 U233 ( .A1(\data_i[29][8] ), .A2(n695), .B1(\data_i[28][8] ), .B2(
        n696), .ZN(n168) );
  AOI22D0 U234 ( .A1(\data_i[31][8] ), .A2(n697), .B1(\data_i[30][8] ), .B2(
        n698), .ZN(n169) );
  ND4D0 U235 ( .A1(n166), .A2(n167), .A3(n168), .A4(n169), .ZN(n170) );
  AOI22D0 U236 ( .A1(\data_i[1][8] ), .A2(n667), .B1(\data_i[0][8] ), .B2(n668), .ZN(n171) );
  AOI22D0 U237 ( .A1(\data_i[3][8] ), .A2(n669), .B1(\data_i[2][8] ), .B2(n670), .ZN(n172) );
  AOI22D0 U238 ( .A1(\data_i[5][8] ), .A2(n671), .B1(\data_i[4][8] ), .B2(n672), .ZN(n173) );
  AOI22D0 U239 ( .A1(\data_i[7][8] ), .A2(n673), .B1(\data_i[6][8] ), .B2(n674), .ZN(n174) );
  ND4D0 U240 ( .A1(n171), .A2(n172), .A3(n173), .A4(n174), .ZN(n175) );
  AOI22D0 U241 ( .A1(\data_i[9][8] ), .A2(n675), .B1(\data_i[8][8] ), .B2(n676), .ZN(n176) );
  AOI22D0 U242 ( .A1(\data_i[11][8] ), .A2(n677), .B1(\data_i[10][8] ), .B2(
        n678), .ZN(n177) );
  AOI22D0 U243 ( .A1(\data_i[13][8] ), .A2(n679), .B1(\data_i[12][8] ), .B2(
        n680), .ZN(n178) );
  AOI22D0 U244 ( .A1(\data_i[15][8] ), .A2(n681), .B1(\data_i[14][8] ), .B2(
        n682), .ZN(n179) );
  ND4D0 U245 ( .A1(n176), .A2(n177), .A3(n178), .A4(n179), .ZN(n180) );
  OR4D0 U246 ( .A1(n165), .A2(n170), .A3(n175), .A4(n180), .Z(data_o[8]) );
  AOI22D0 U247 ( .A1(\data_i[17][9] ), .A2(n683), .B1(\data_i[16][9] ), .B2(
        n684), .ZN(n181) );
  AOI22D0 U248 ( .A1(\data_i[19][9] ), .A2(n685), .B1(\data_i[18][9] ), .B2(
        n686), .ZN(n182) );
  AOI22D0 U249 ( .A1(\data_i[21][9] ), .A2(n687), .B1(\data_i[20][9] ), .B2(
        n688), .ZN(n183) );
  AOI22D0 U250 ( .A1(\data_i[23][9] ), .A2(n689), .B1(\data_i[22][9] ), .B2(
        n690), .ZN(n184) );
  ND4D0 U251 ( .A1(n181), .A2(n182), .A3(n183), .A4(n184), .ZN(n185) );
  AOI22D0 U252 ( .A1(\data_i[25][9] ), .A2(n691), .B1(\data_i[24][9] ), .B2(
        n692), .ZN(n186) );
  AOI22D0 U253 ( .A1(\data_i[27][9] ), .A2(n693), .B1(\data_i[26][9] ), .B2(
        n694), .ZN(n187) );
  AOI22D0 U254 ( .A1(\data_i[29][9] ), .A2(n695), .B1(\data_i[28][9] ), .B2(
        n696), .ZN(n188) );
  AOI22D0 U255 ( .A1(\data_i[31][9] ), .A2(n697), .B1(\data_i[30][9] ), .B2(
        n698), .ZN(n189) );
  ND4D0 U256 ( .A1(n186), .A2(n187), .A3(n188), .A4(n189), .ZN(n190) );
  AOI22D0 U257 ( .A1(\data_i[1][9] ), .A2(n667), .B1(\data_i[0][9] ), .B2(n668), .ZN(n191) );
  AOI22D0 U258 ( .A1(\data_i[3][9] ), .A2(n669), .B1(\data_i[2][9] ), .B2(n670), .ZN(n192) );
  AOI22D0 U259 ( .A1(\data_i[5][9] ), .A2(n671), .B1(\data_i[4][9] ), .B2(n672), .ZN(n193) );
  AOI22D0 U260 ( .A1(\data_i[7][9] ), .A2(n673), .B1(\data_i[6][9] ), .B2(n674), .ZN(n194) );
  ND4D0 U261 ( .A1(n191), .A2(n192), .A3(n193), .A4(n194), .ZN(n195) );
  AOI22D0 U262 ( .A1(\data_i[9][9] ), .A2(n675), .B1(\data_i[8][9] ), .B2(n676), .ZN(n196) );
  AOI22D0 U263 ( .A1(\data_i[11][9] ), .A2(n677), .B1(\data_i[10][9] ), .B2(
        n678), .ZN(n197) );
  AOI22D0 U264 ( .A1(\data_i[13][9] ), .A2(n679), .B1(\data_i[12][9] ), .B2(
        n680), .ZN(n198) );
  AOI22D0 U265 ( .A1(\data_i[15][9] ), .A2(n681), .B1(\data_i[14][9] ), .B2(
        n682), .ZN(n199) );
  ND4D0 U266 ( .A1(n196), .A2(n197), .A3(n198), .A4(n199), .ZN(n200) );
  OR4D0 U267 ( .A1(n185), .A2(n190), .A3(n195), .A4(n200), .Z(data_o[9]) );
  AOI22D0 U268 ( .A1(\data_i[17][10] ), .A2(n683), .B1(\data_i[16][10] ), .B2(
        n684), .ZN(n201) );
  AOI22D0 U269 ( .A1(\data_i[19][10] ), .A2(n685), .B1(\data_i[18][10] ), .B2(
        n686), .ZN(n202) );
  AOI22D0 U270 ( .A1(\data_i[21][10] ), .A2(n687), .B1(\data_i[20][10] ), .B2(
        n688), .ZN(n203) );
  AOI22D0 U271 ( .A1(\data_i[23][10] ), .A2(n689), .B1(\data_i[22][10] ), .B2(
        n690), .ZN(n204) );
  ND4D0 U272 ( .A1(n201), .A2(n202), .A3(n203), .A4(n204), .ZN(n205) );
  AOI22D0 U273 ( .A1(\data_i[25][10] ), .A2(n691), .B1(\data_i[24][10] ), .B2(
        n692), .ZN(n206) );
  AOI22D0 U274 ( .A1(\data_i[27][10] ), .A2(n693), .B1(\data_i[26][10] ), .B2(
        n694), .ZN(n207) );
  AOI22D0 U275 ( .A1(\data_i[29][10] ), .A2(n695), .B1(\data_i[28][10] ), .B2(
        n696), .ZN(n208) );
  AOI22D0 U276 ( .A1(\data_i[31][10] ), .A2(n697), .B1(\data_i[30][10] ), .B2(
        n698), .ZN(n209) );
  ND4D0 U277 ( .A1(n206), .A2(n207), .A3(n208), .A4(n209), .ZN(n210) );
  AOI22D0 U278 ( .A1(\data_i[1][10] ), .A2(n667), .B1(\data_i[0][10] ), .B2(
        n668), .ZN(n211) );
  AOI22D0 U279 ( .A1(\data_i[3][10] ), .A2(n669), .B1(\data_i[2][10] ), .B2(
        n670), .ZN(n212) );
  AOI22D0 U280 ( .A1(\data_i[5][10] ), .A2(n671), .B1(\data_i[4][10] ), .B2(
        n672), .ZN(n213) );
  AOI22D0 U281 ( .A1(\data_i[7][10] ), .A2(n673), .B1(\data_i[6][10] ), .B2(
        n674), .ZN(n214) );
  ND4D0 U282 ( .A1(n211), .A2(n212), .A3(n213), .A4(n214), .ZN(n215) );
  AOI22D0 U283 ( .A1(\data_i[9][10] ), .A2(n675), .B1(\data_i[8][10] ), .B2(
        n676), .ZN(n216) );
  AOI22D0 U284 ( .A1(\data_i[11][10] ), .A2(n677), .B1(\data_i[10][10] ), .B2(
        n678), .ZN(n217) );
  AOI22D0 U285 ( .A1(\data_i[13][10] ), .A2(n679), .B1(\data_i[12][10] ), .B2(
        n680), .ZN(n218) );
  AOI22D0 U286 ( .A1(\data_i[15][10] ), .A2(n681), .B1(\data_i[14][10] ), .B2(
        n682), .ZN(n219) );
  ND4D0 U287 ( .A1(n216), .A2(n217), .A3(n218), .A4(n219), .ZN(n220) );
  OR4D0 U288 ( .A1(n205), .A2(n210), .A3(n215), .A4(n220), .Z(data_o[10]) );
  AOI22D0 U289 ( .A1(\data_i[17][11] ), .A2(n683), .B1(\data_i[16][11] ), .B2(
        n684), .ZN(n221) );
  AOI22D0 U290 ( .A1(\data_i[19][11] ), .A2(n685), .B1(\data_i[18][11] ), .B2(
        n686), .ZN(n222) );
  AOI22D0 U291 ( .A1(\data_i[21][11] ), .A2(n687), .B1(\data_i[20][11] ), .B2(
        n688), .ZN(n223) );
  AOI22D0 U292 ( .A1(\data_i[23][11] ), .A2(n689), .B1(\data_i[22][11] ), .B2(
        n690), .ZN(n224) );
  ND4D0 U293 ( .A1(n221), .A2(n222), .A3(n223), .A4(n224), .ZN(n225) );
  AOI22D0 U294 ( .A1(\data_i[25][11] ), .A2(n691), .B1(\data_i[24][11] ), .B2(
        n692), .ZN(n226) );
  AOI22D0 U295 ( .A1(\data_i[27][11] ), .A2(n693), .B1(\data_i[26][11] ), .B2(
        n694), .ZN(n227) );
  AOI22D0 U296 ( .A1(\data_i[29][11] ), .A2(n695), .B1(\data_i[28][11] ), .B2(
        n696), .ZN(n228) );
  AOI22D0 U297 ( .A1(\data_i[31][11] ), .A2(n697), .B1(\data_i[30][11] ), .B2(
        n698), .ZN(n229) );
  ND4D0 U298 ( .A1(n226), .A2(n227), .A3(n228), .A4(n229), .ZN(n230) );
  AOI22D0 U299 ( .A1(\data_i[1][11] ), .A2(n667), .B1(\data_i[0][11] ), .B2(
        n668), .ZN(n231) );
  AOI22D0 U300 ( .A1(\data_i[3][11] ), .A2(n669), .B1(\data_i[2][11] ), .B2(
        n670), .ZN(n232) );
  AOI22D0 U301 ( .A1(\data_i[5][11] ), .A2(n671), .B1(\data_i[4][11] ), .B2(
        n672), .ZN(n233) );
  AOI22D0 U302 ( .A1(\data_i[7][11] ), .A2(n673), .B1(\data_i[6][11] ), .B2(
        n674), .ZN(n234) );
  ND4D0 U303 ( .A1(n231), .A2(n232), .A3(n233), .A4(n234), .ZN(n235) );
  AOI22D0 U304 ( .A1(\data_i[9][11] ), .A2(n675), .B1(\data_i[8][11] ), .B2(
        n676), .ZN(n236) );
  AOI22D0 U305 ( .A1(\data_i[11][11] ), .A2(n677), .B1(\data_i[10][11] ), .B2(
        n678), .ZN(n237) );
  AOI22D0 U306 ( .A1(\data_i[13][11] ), .A2(n679), .B1(\data_i[12][11] ), .B2(
        n680), .ZN(n238) );
  AOI22D0 U307 ( .A1(\data_i[15][11] ), .A2(n681), .B1(\data_i[14][11] ), .B2(
        n682), .ZN(n239) );
  ND4D0 U308 ( .A1(n236), .A2(n237), .A3(n238), .A4(n239), .ZN(n240) );
  OR4D0 U309 ( .A1(n225), .A2(n230), .A3(n235), .A4(n240), .Z(data_o[11]) );
  AOI22D0 U310 ( .A1(\data_i[17][12] ), .A2(n683), .B1(\data_i[16][12] ), .B2(
        n684), .ZN(n241) );
  AOI22D0 U311 ( .A1(\data_i[19][12] ), .A2(n685), .B1(\data_i[18][12] ), .B2(
        n686), .ZN(n242) );
  AOI22D0 U312 ( .A1(\data_i[21][12] ), .A2(n687), .B1(\data_i[20][12] ), .B2(
        n688), .ZN(n243) );
  AOI22D0 U313 ( .A1(\data_i[23][12] ), .A2(n689), .B1(\data_i[22][12] ), .B2(
        n690), .ZN(n244) );
  ND4D0 U314 ( .A1(n241), .A2(n242), .A3(n243), .A4(n244), .ZN(n245) );
  AOI22D0 U315 ( .A1(\data_i[25][12] ), .A2(n691), .B1(\data_i[24][12] ), .B2(
        n692), .ZN(n246) );
  AOI22D0 U316 ( .A1(\data_i[27][12] ), .A2(n693), .B1(\data_i[26][12] ), .B2(
        n694), .ZN(n247) );
  AOI22D0 U317 ( .A1(\data_i[29][12] ), .A2(n695), .B1(\data_i[28][12] ), .B2(
        n696), .ZN(n248) );
  AOI22D0 U318 ( .A1(\data_i[31][12] ), .A2(n697), .B1(\data_i[30][12] ), .B2(
        n698), .ZN(n249) );
  ND4D0 U319 ( .A1(n246), .A2(n247), .A3(n248), .A4(n249), .ZN(n250) );
  AOI22D0 U320 ( .A1(\data_i[1][12] ), .A2(n667), .B1(\data_i[0][12] ), .B2(
        n668), .ZN(n251) );
  AOI22D0 U321 ( .A1(\data_i[3][12] ), .A2(n669), .B1(\data_i[2][12] ), .B2(
        n670), .ZN(n252) );
  AOI22D0 U322 ( .A1(\data_i[5][12] ), .A2(n671), .B1(\data_i[4][12] ), .B2(
        n672), .ZN(n253) );
  AOI22D0 U323 ( .A1(\data_i[7][12] ), .A2(n673), .B1(\data_i[6][12] ), .B2(
        n674), .ZN(n254) );
  ND4D0 U324 ( .A1(n251), .A2(n252), .A3(n253), .A4(n254), .ZN(n255) );
  AOI22D0 U325 ( .A1(\data_i[9][12] ), .A2(n675), .B1(\data_i[8][12] ), .B2(
        n676), .ZN(n256) );
  AOI22D0 U326 ( .A1(\data_i[11][12] ), .A2(n677), .B1(\data_i[10][12] ), .B2(
        n678), .ZN(n257) );
  AOI22D0 U327 ( .A1(\data_i[13][12] ), .A2(n679), .B1(\data_i[12][12] ), .B2(
        n680), .ZN(n258) );
  AOI22D0 U328 ( .A1(\data_i[15][12] ), .A2(n681), .B1(\data_i[14][12] ), .B2(
        n682), .ZN(n259) );
  ND4D0 U329 ( .A1(n256), .A2(n257), .A3(n258), .A4(n259), .ZN(n260) );
  OR4D0 U330 ( .A1(n245), .A2(n250), .A3(n255), .A4(n260), .Z(data_o[12]) );
  AOI22D0 U331 ( .A1(\data_i[17][13] ), .A2(n683), .B1(\data_i[16][13] ), .B2(
        n684), .ZN(n261) );
  AOI22D0 U332 ( .A1(\data_i[19][13] ), .A2(n685), .B1(\data_i[18][13] ), .B2(
        n686), .ZN(n262) );
  AOI22D0 U333 ( .A1(\data_i[21][13] ), .A2(n687), .B1(\data_i[20][13] ), .B2(
        n688), .ZN(n263) );
  AOI22D0 U334 ( .A1(\data_i[23][13] ), .A2(n689), .B1(\data_i[22][13] ), .B2(
        n690), .ZN(n264) );
  ND4D0 U335 ( .A1(n261), .A2(n262), .A3(n263), .A4(n264), .ZN(n265) );
  AOI22D0 U336 ( .A1(\data_i[25][13] ), .A2(n691), .B1(\data_i[24][13] ), .B2(
        n692), .ZN(n266) );
  AOI22D0 U337 ( .A1(\data_i[27][13] ), .A2(n693), .B1(\data_i[26][13] ), .B2(
        n694), .ZN(n267) );
  AOI22D0 U338 ( .A1(\data_i[29][13] ), .A2(n695), .B1(\data_i[28][13] ), .B2(
        n696), .ZN(n268) );
  AOI22D0 U339 ( .A1(\data_i[31][13] ), .A2(n697), .B1(\data_i[30][13] ), .B2(
        n698), .ZN(n269) );
  ND4D0 U340 ( .A1(n266), .A2(n267), .A3(n268), .A4(n269), .ZN(n270) );
  AOI22D0 U341 ( .A1(\data_i[1][13] ), .A2(n667), .B1(\data_i[0][13] ), .B2(
        n668), .ZN(n271) );
  AOI22D0 U342 ( .A1(\data_i[3][13] ), .A2(n669), .B1(\data_i[2][13] ), .B2(
        n670), .ZN(n272) );
  AOI22D0 U343 ( .A1(\data_i[5][13] ), .A2(n671), .B1(\data_i[4][13] ), .B2(
        n672), .ZN(n273) );
  AOI22D0 U344 ( .A1(\data_i[7][13] ), .A2(n673), .B1(\data_i[6][13] ), .B2(
        n674), .ZN(n274) );
  ND4D0 U345 ( .A1(n271), .A2(n272), .A3(n273), .A4(n274), .ZN(n275) );
  AOI22D0 U346 ( .A1(\data_i[9][13] ), .A2(n675), .B1(\data_i[8][13] ), .B2(
        n676), .ZN(n276) );
  AOI22D0 U347 ( .A1(\data_i[11][13] ), .A2(n677), .B1(\data_i[10][13] ), .B2(
        n678), .ZN(n277) );
  AOI22D0 U348 ( .A1(\data_i[13][13] ), .A2(n679), .B1(\data_i[12][13] ), .B2(
        n680), .ZN(n278) );
  AOI22D0 U349 ( .A1(\data_i[15][13] ), .A2(n681), .B1(\data_i[14][13] ), .B2(
        n682), .ZN(n279) );
  ND4D0 U350 ( .A1(n276), .A2(n277), .A3(n278), .A4(n279), .ZN(n280) );
  OR4D0 U351 ( .A1(n265), .A2(n270), .A3(n275), .A4(n280), .Z(data_o[13]) );
  AOI22D0 U352 ( .A1(\data_i[17][14] ), .A2(n683), .B1(\data_i[16][14] ), .B2(
        n684), .ZN(n281) );
  AOI22D0 U353 ( .A1(\data_i[19][14] ), .A2(n685), .B1(\data_i[18][14] ), .B2(
        n686), .ZN(n282) );
  AOI22D0 U354 ( .A1(\data_i[21][14] ), .A2(n687), .B1(\data_i[20][14] ), .B2(
        n688), .ZN(n283) );
  AOI22D0 U355 ( .A1(\data_i[23][14] ), .A2(n689), .B1(\data_i[22][14] ), .B2(
        n690), .ZN(n284) );
  ND4D0 U356 ( .A1(n281), .A2(n282), .A3(n283), .A4(n284), .ZN(n285) );
  AOI22D0 U357 ( .A1(\data_i[25][14] ), .A2(n691), .B1(\data_i[24][14] ), .B2(
        n692), .ZN(n286) );
  AOI22D0 U358 ( .A1(\data_i[27][14] ), .A2(n693), .B1(\data_i[26][14] ), .B2(
        n694), .ZN(n287) );
  AOI22D0 U359 ( .A1(\data_i[29][14] ), .A2(n695), .B1(\data_i[28][14] ), .B2(
        n696), .ZN(n288) );
  AOI22D0 U360 ( .A1(\data_i[31][14] ), .A2(n697), .B1(\data_i[30][14] ), .B2(
        n698), .ZN(n289) );
  ND4D0 U361 ( .A1(n286), .A2(n287), .A3(n288), .A4(n289), .ZN(n290) );
  AOI22D0 U362 ( .A1(\data_i[1][14] ), .A2(n667), .B1(\data_i[0][14] ), .B2(
        n668), .ZN(n291) );
  AOI22D0 U363 ( .A1(\data_i[3][14] ), .A2(n669), .B1(\data_i[2][14] ), .B2(
        n670), .ZN(n292) );
  AOI22D0 U364 ( .A1(\data_i[5][14] ), .A2(n671), .B1(\data_i[4][14] ), .B2(
        n672), .ZN(n293) );
  AOI22D0 U365 ( .A1(\data_i[7][14] ), .A2(n673), .B1(\data_i[6][14] ), .B2(
        n674), .ZN(n294) );
  ND4D0 U366 ( .A1(n291), .A2(n292), .A3(n293), .A4(n294), .ZN(n295) );
  AOI22D0 U367 ( .A1(\data_i[9][14] ), .A2(n675), .B1(\data_i[8][14] ), .B2(
        n676), .ZN(n296) );
  AOI22D0 U368 ( .A1(\data_i[11][14] ), .A2(n677), .B1(\data_i[10][14] ), .B2(
        n678), .ZN(n297) );
  AOI22D0 U369 ( .A1(\data_i[13][14] ), .A2(n679), .B1(\data_i[12][14] ), .B2(
        n680), .ZN(n298) );
  AOI22D0 U370 ( .A1(\data_i[15][14] ), .A2(n681), .B1(\data_i[14][14] ), .B2(
        n682), .ZN(n299) );
  ND4D0 U371 ( .A1(n296), .A2(n297), .A3(n298), .A4(n299), .ZN(n300) );
  OR4D0 U372 ( .A1(n285), .A2(n290), .A3(n295), .A4(n300), .Z(data_o[14]) );
  AOI22D0 U373 ( .A1(\data_i[17][15] ), .A2(n683), .B1(\data_i[16][15] ), .B2(
        n684), .ZN(n301) );
  AOI22D0 U374 ( .A1(\data_i[19][15] ), .A2(n685), .B1(\data_i[18][15] ), .B2(
        n686), .ZN(n302) );
  AOI22D0 U375 ( .A1(\data_i[21][15] ), .A2(n687), .B1(\data_i[20][15] ), .B2(
        n688), .ZN(n303) );
  AOI22D0 U376 ( .A1(\data_i[23][15] ), .A2(n689), .B1(\data_i[22][15] ), .B2(
        n690), .ZN(n304) );
  ND4D0 U377 ( .A1(n301), .A2(n302), .A3(n303), .A4(n304), .ZN(n305) );
  AOI22D0 U378 ( .A1(\data_i[25][15] ), .A2(n691), .B1(\data_i[24][15] ), .B2(
        n692), .ZN(n306) );
  AOI22D0 U379 ( .A1(\data_i[27][15] ), .A2(n693), .B1(\data_i[26][15] ), .B2(
        n694), .ZN(n307) );
  AOI22D0 U380 ( .A1(\data_i[29][15] ), .A2(n695), .B1(\data_i[28][15] ), .B2(
        n696), .ZN(n308) );
  AOI22D0 U381 ( .A1(\data_i[31][15] ), .A2(n697), .B1(\data_i[30][15] ), .B2(
        n698), .ZN(n309) );
  ND4D0 U382 ( .A1(n306), .A2(n307), .A3(n308), .A4(n309), .ZN(n310) );
  AOI22D0 U383 ( .A1(\data_i[1][15] ), .A2(n667), .B1(\data_i[0][15] ), .B2(
        n668), .ZN(n311) );
  AOI22D0 U384 ( .A1(\data_i[3][15] ), .A2(n669), .B1(\data_i[2][15] ), .B2(
        n670), .ZN(n312) );
  AOI22D0 U385 ( .A1(\data_i[5][15] ), .A2(n671), .B1(\data_i[4][15] ), .B2(
        n672), .ZN(n313) );
  AOI22D0 U386 ( .A1(\data_i[7][15] ), .A2(n673), .B1(\data_i[6][15] ), .B2(
        n674), .ZN(n314) );
  ND4D0 U387 ( .A1(n311), .A2(n312), .A3(n313), .A4(n314), .ZN(n315) );
  AOI22D0 U388 ( .A1(\data_i[9][15] ), .A2(n675), .B1(\data_i[8][15] ), .B2(
        n676), .ZN(n316) );
  AOI22D0 U389 ( .A1(\data_i[11][15] ), .A2(n677), .B1(\data_i[10][15] ), .B2(
        n678), .ZN(n317) );
  AOI22D0 U390 ( .A1(\data_i[13][15] ), .A2(n679), .B1(\data_i[12][15] ), .B2(
        n680), .ZN(n318) );
  AOI22D0 U391 ( .A1(\data_i[15][15] ), .A2(n681), .B1(\data_i[14][15] ), .B2(
        n682), .ZN(n319) );
  ND4D0 U392 ( .A1(n316), .A2(n317), .A3(n318), .A4(n319), .ZN(n320) );
  OR4D0 U393 ( .A1(n305), .A2(n310), .A3(n315), .A4(n320), .Z(data_o[15]) );
  AOI22D0 U394 ( .A1(\data_i[17][16] ), .A2(n683), .B1(\data_i[16][16] ), .B2(
        n684), .ZN(n321) );
  AOI22D0 U395 ( .A1(\data_i[19][16] ), .A2(n685), .B1(\data_i[18][16] ), .B2(
        n686), .ZN(n322) );
  AOI22D0 U396 ( .A1(\data_i[21][16] ), .A2(n687), .B1(\data_i[20][16] ), .B2(
        n688), .ZN(n323) );
  AOI22D0 U397 ( .A1(\data_i[23][16] ), .A2(n689), .B1(\data_i[22][16] ), .B2(
        n690), .ZN(n324) );
  ND4D0 U398 ( .A1(n321), .A2(n322), .A3(n323), .A4(n324), .ZN(n325) );
  AOI22D0 U399 ( .A1(\data_i[25][16] ), .A2(n691), .B1(\data_i[24][16] ), .B2(
        n692), .ZN(n326) );
  AOI22D0 U400 ( .A1(\data_i[27][16] ), .A2(n693), .B1(\data_i[26][16] ), .B2(
        n694), .ZN(n327) );
  AOI22D0 U401 ( .A1(\data_i[29][16] ), .A2(n695), .B1(\data_i[28][16] ), .B2(
        n696), .ZN(n328) );
  AOI22D0 U402 ( .A1(\data_i[31][16] ), .A2(n697), .B1(\data_i[30][16] ), .B2(
        n698), .ZN(n329) );
  ND4D0 U403 ( .A1(n326), .A2(n327), .A3(n328), .A4(n329), .ZN(n330) );
  AOI22D0 U404 ( .A1(\data_i[1][16] ), .A2(n667), .B1(\data_i[0][16] ), .B2(
        n668), .ZN(n331) );
  AOI22D0 U405 ( .A1(\data_i[3][16] ), .A2(n669), .B1(\data_i[2][16] ), .B2(
        n670), .ZN(n332) );
  AOI22D0 U406 ( .A1(\data_i[5][16] ), .A2(n671), .B1(\data_i[4][16] ), .B2(
        n672), .ZN(n333) );
  AOI22D0 U407 ( .A1(\data_i[7][16] ), .A2(n673), .B1(\data_i[6][16] ), .B2(
        n674), .ZN(n334) );
  ND4D0 U408 ( .A1(n331), .A2(n332), .A3(n333), .A4(n334), .ZN(n335) );
  AOI22D0 U409 ( .A1(\data_i[9][16] ), .A2(n675), .B1(\data_i[8][16] ), .B2(
        n676), .ZN(n336) );
  AOI22D0 U410 ( .A1(\data_i[11][16] ), .A2(n677), .B1(\data_i[10][16] ), .B2(
        n678), .ZN(n337) );
  AOI22D0 U411 ( .A1(\data_i[13][16] ), .A2(n679), .B1(\data_i[12][16] ), .B2(
        n680), .ZN(n338) );
  AOI22D0 U412 ( .A1(\data_i[15][16] ), .A2(n681), .B1(\data_i[14][16] ), .B2(
        n682), .ZN(n339) );
  ND4D0 U413 ( .A1(n336), .A2(n337), .A3(n338), .A4(n339), .ZN(n340) );
  OR4D0 U414 ( .A1(n325), .A2(n330), .A3(n335), .A4(n340), .Z(data_o[16]) );
  AOI22D0 U415 ( .A1(\data_i[17][17] ), .A2(n683), .B1(\data_i[16][17] ), .B2(
        n684), .ZN(n341) );
  AOI22D0 U416 ( .A1(\data_i[19][17] ), .A2(n685), .B1(\data_i[18][17] ), .B2(
        n686), .ZN(n342) );
  AOI22D0 U417 ( .A1(\data_i[21][17] ), .A2(n687), .B1(\data_i[20][17] ), .B2(
        n688), .ZN(n343) );
  AOI22D0 U418 ( .A1(\data_i[23][17] ), .A2(n689), .B1(\data_i[22][17] ), .B2(
        n690), .ZN(n344) );
  ND4D0 U419 ( .A1(n341), .A2(n342), .A3(n343), .A4(n344), .ZN(n345) );
  AOI22D0 U420 ( .A1(\data_i[25][17] ), .A2(n691), .B1(\data_i[24][17] ), .B2(
        n692), .ZN(n346) );
  AOI22D0 U421 ( .A1(\data_i[27][17] ), .A2(n693), .B1(\data_i[26][17] ), .B2(
        n694), .ZN(n347) );
  AOI22D0 U422 ( .A1(\data_i[29][17] ), .A2(n695), .B1(\data_i[28][17] ), .B2(
        n696), .ZN(n348) );
  AOI22D0 U423 ( .A1(\data_i[31][17] ), .A2(n697), .B1(\data_i[30][17] ), .B2(
        n698), .ZN(n349) );
  ND4D0 U424 ( .A1(n346), .A2(n347), .A3(n348), .A4(n349), .ZN(n350) );
  AOI22D0 U425 ( .A1(\data_i[1][17] ), .A2(n667), .B1(\data_i[0][17] ), .B2(
        n668), .ZN(n351) );
  AOI22D0 U426 ( .A1(\data_i[3][17] ), .A2(n669), .B1(\data_i[2][17] ), .B2(
        n670), .ZN(n352) );
  AOI22D0 U427 ( .A1(\data_i[5][17] ), .A2(n671), .B1(\data_i[4][17] ), .B2(
        n672), .ZN(n353) );
  AOI22D0 U428 ( .A1(\data_i[7][17] ), .A2(n673), .B1(\data_i[6][17] ), .B2(
        n674), .ZN(n354) );
  ND4D0 U429 ( .A1(n351), .A2(n352), .A3(n353), .A4(n354), .ZN(n355) );
  AOI22D0 U430 ( .A1(\data_i[9][17] ), .A2(n675), .B1(\data_i[8][17] ), .B2(
        n676), .ZN(n356) );
  AOI22D0 U431 ( .A1(\data_i[11][17] ), .A2(n677), .B1(\data_i[10][17] ), .B2(
        n678), .ZN(n357) );
  AOI22D0 U432 ( .A1(\data_i[13][17] ), .A2(n679), .B1(\data_i[12][17] ), .B2(
        n680), .ZN(n358) );
  AOI22D0 U433 ( .A1(\data_i[15][17] ), .A2(n681), .B1(\data_i[14][17] ), .B2(
        n682), .ZN(n359) );
  ND4D0 U434 ( .A1(n356), .A2(n357), .A3(n358), .A4(n359), .ZN(n360) );
  OR4D0 U435 ( .A1(n345), .A2(n350), .A3(n355), .A4(n360), .Z(data_o[17]) );
  AOI22D0 U436 ( .A1(\data_i[17][18] ), .A2(n683), .B1(\data_i[16][18] ), .B2(
        n684), .ZN(n361) );
  AOI22D0 U437 ( .A1(\data_i[19][18] ), .A2(n685), .B1(\data_i[18][18] ), .B2(
        n686), .ZN(n362) );
  AOI22D0 U438 ( .A1(\data_i[21][18] ), .A2(n687), .B1(\data_i[20][18] ), .B2(
        n688), .ZN(n363) );
  AOI22D0 U439 ( .A1(\data_i[23][18] ), .A2(n689), .B1(\data_i[22][18] ), .B2(
        n690), .ZN(n364) );
  ND4D0 U440 ( .A1(n361), .A2(n362), .A3(n363), .A4(n364), .ZN(n365) );
  AOI22D0 U441 ( .A1(\data_i[25][18] ), .A2(n691), .B1(\data_i[24][18] ), .B2(
        n692), .ZN(n366) );
  AOI22D0 U442 ( .A1(\data_i[27][18] ), .A2(n693), .B1(\data_i[26][18] ), .B2(
        n694), .ZN(n367) );
  AOI22D0 U443 ( .A1(\data_i[29][18] ), .A2(n695), .B1(\data_i[28][18] ), .B2(
        n696), .ZN(n368) );
  AOI22D0 U444 ( .A1(\data_i[31][18] ), .A2(n697), .B1(\data_i[30][18] ), .B2(
        n698), .ZN(n369) );
  ND4D0 U445 ( .A1(n366), .A2(n367), .A3(n368), .A4(n369), .ZN(n370) );
  AOI22D0 U446 ( .A1(\data_i[1][18] ), .A2(n667), .B1(\data_i[0][18] ), .B2(
        n668), .ZN(n371) );
  AOI22D0 U447 ( .A1(\data_i[3][18] ), .A2(n669), .B1(\data_i[2][18] ), .B2(
        n670), .ZN(n372) );
  AOI22D0 U448 ( .A1(\data_i[5][18] ), .A2(n671), .B1(\data_i[4][18] ), .B2(
        n672), .ZN(n373) );
  AOI22D0 U449 ( .A1(\data_i[7][18] ), .A2(n673), .B1(\data_i[6][18] ), .B2(
        n674), .ZN(n374) );
  ND4D0 U450 ( .A1(n371), .A2(n372), .A3(n373), .A4(n374), .ZN(n375) );
  AOI22D0 U451 ( .A1(\data_i[9][18] ), .A2(n675), .B1(\data_i[8][18] ), .B2(
        n676), .ZN(n376) );
  AOI22D0 U452 ( .A1(\data_i[11][18] ), .A2(n677), .B1(\data_i[10][18] ), .B2(
        n678), .ZN(n377) );
  AOI22D0 U453 ( .A1(\data_i[13][18] ), .A2(n679), .B1(\data_i[12][18] ), .B2(
        n680), .ZN(n378) );
  AOI22D0 U454 ( .A1(\data_i[15][18] ), .A2(n681), .B1(\data_i[14][18] ), .B2(
        n682), .ZN(n379) );
  ND4D0 U455 ( .A1(n376), .A2(n377), .A3(n378), .A4(n379), .ZN(n380) );
  OR4D0 U456 ( .A1(n365), .A2(n370), .A3(n375), .A4(n380), .Z(data_o[18]) );
  AOI22D0 U457 ( .A1(\data_i[17][19] ), .A2(n683), .B1(\data_i[16][19] ), .B2(
        n684), .ZN(n381) );
  AOI22D0 U458 ( .A1(\data_i[19][19] ), .A2(n685), .B1(\data_i[18][19] ), .B2(
        n686), .ZN(n382) );
  AOI22D0 U459 ( .A1(\data_i[21][19] ), .A2(n687), .B1(\data_i[20][19] ), .B2(
        n688), .ZN(n383) );
  AOI22D0 U460 ( .A1(\data_i[23][19] ), .A2(n689), .B1(\data_i[22][19] ), .B2(
        n690), .ZN(n384) );
  ND4D0 U461 ( .A1(n381), .A2(n382), .A3(n383), .A4(n384), .ZN(n385) );
  AOI22D0 U462 ( .A1(\data_i[25][19] ), .A2(n691), .B1(\data_i[24][19] ), .B2(
        n692), .ZN(n386) );
  AOI22D0 U463 ( .A1(\data_i[27][19] ), .A2(n693), .B1(\data_i[26][19] ), .B2(
        n694), .ZN(n387) );
  AOI22D0 U464 ( .A1(\data_i[29][19] ), .A2(n695), .B1(\data_i[28][19] ), .B2(
        n696), .ZN(n388) );
  AOI22D0 U465 ( .A1(\data_i[31][19] ), .A2(n697), .B1(\data_i[30][19] ), .B2(
        n698), .ZN(n389) );
  ND4D0 U466 ( .A1(n386), .A2(n387), .A3(n388), .A4(n389), .ZN(n390) );
  AOI22D0 U467 ( .A1(\data_i[1][19] ), .A2(n667), .B1(\data_i[0][19] ), .B2(
        n668), .ZN(n391) );
  AOI22D0 U468 ( .A1(\data_i[3][19] ), .A2(n669), .B1(\data_i[2][19] ), .B2(
        n670), .ZN(n392) );
  AOI22D0 U469 ( .A1(\data_i[5][19] ), .A2(n671), .B1(\data_i[4][19] ), .B2(
        n672), .ZN(n393) );
  AOI22D0 U470 ( .A1(\data_i[7][19] ), .A2(n673), .B1(\data_i[6][19] ), .B2(
        n674), .ZN(n394) );
  ND4D0 U471 ( .A1(n391), .A2(n392), .A3(n393), .A4(n394), .ZN(n395) );
  AOI22D0 U472 ( .A1(\data_i[9][19] ), .A2(n675), .B1(\data_i[8][19] ), .B2(
        n676), .ZN(n396) );
  AOI22D0 U473 ( .A1(\data_i[11][19] ), .A2(n677), .B1(\data_i[10][19] ), .B2(
        n678), .ZN(n397) );
  AOI22D0 U474 ( .A1(\data_i[13][19] ), .A2(n679), .B1(\data_i[12][19] ), .B2(
        n680), .ZN(n398) );
  AOI22D0 U475 ( .A1(\data_i[15][19] ), .A2(n681), .B1(\data_i[14][19] ), .B2(
        n682), .ZN(n399) );
  ND4D0 U476 ( .A1(n396), .A2(n397), .A3(n398), .A4(n399), .ZN(n400) );
  OR4D0 U477 ( .A1(n385), .A2(n390), .A3(n395), .A4(n400), .Z(data_o[19]) );
  AOI22D0 U478 ( .A1(\data_i[17][20] ), .A2(n683), .B1(\data_i[16][20] ), .B2(
        n684), .ZN(n401) );
  AOI22D0 U479 ( .A1(\data_i[19][20] ), .A2(n685), .B1(\data_i[18][20] ), .B2(
        n686), .ZN(n402) );
  AOI22D0 U480 ( .A1(\data_i[21][20] ), .A2(n687), .B1(\data_i[20][20] ), .B2(
        n688), .ZN(n403) );
  AOI22D0 U481 ( .A1(\data_i[23][20] ), .A2(n689), .B1(\data_i[22][20] ), .B2(
        n690), .ZN(n404) );
  ND4D0 U482 ( .A1(n401), .A2(n402), .A3(n403), .A4(n404), .ZN(n405) );
  AOI22D0 U483 ( .A1(\data_i[25][20] ), .A2(n691), .B1(\data_i[24][20] ), .B2(
        n692), .ZN(n406) );
  AOI22D0 U484 ( .A1(\data_i[27][20] ), .A2(n693), .B1(\data_i[26][20] ), .B2(
        n694), .ZN(n407) );
  AOI22D0 U485 ( .A1(\data_i[29][20] ), .A2(n695), .B1(\data_i[28][20] ), .B2(
        n696), .ZN(n408) );
  AOI22D0 U486 ( .A1(\data_i[31][20] ), .A2(n697), .B1(\data_i[30][20] ), .B2(
        n698), .ZN(n409) );
  ND4D0 U487 ( .A1(n406), .A2(n407), .A3(n408), .A4(n409), .ZN(n410) );
  AOI22D0 U488 ( .A1(\data_i[1][20] ), .A2(n667), .B1(\data_i[0][20] ), .B2(
        n668), .ZN(n411) );
  AOI22D0 U489 ( .A1(\data_i[3][20] ), .A2(n669), .B1(\data_i[2][20] ), .B2(
        n670), .ZN(n412) );
  AOI22D0 U490 ( .A1(\data_i[5][20] ), .A2(n671), .B1(\data_i[4][20] ), .B2(
        n672), .ZN(n413) );
  AOI22D0 U491 ( .A1(\data_i[7][20] ), .A2(n673), .B1(\data_i[6][20] ), .B2(
        n674), .ZN(n414) );
  ND4D0 U492 ( .A1(n411), .A2(n412), .A3(n413), .A4(n414), .ZN(n415) );
  AOI22D0 U493 ( .A1(\data_i[9][20] ), .A2(n675), .B1(\data_i[8][20] ), .B2(
        n676), .ZN(n416) );
  AOI22D0 U494 ( .A1(\data_i[11][20] ), .A2(n677), .B1(\data_i[10][20] ), .B2(
        n678), .ZN(n417) );
  AOI22D0 U495 ( .A1(\data_i[13][20] ), .A2(n679), .B1(\data_i[12][20] ), .B2(
        n680), .ZN(n418) );
  AOI22D0 U496 ( .A1(\data_i[15][20] ), .A2(n681), .B1(\data_i[14][20] ), .B2(
        n682), .ZN(n419) );
  ND4D0 U497 ( .A1(n416), .A2(n417), .A3(n418), .A4(n419), .ZN(n420) );
  OR4D0 U498 ( .A1(n405), .A2(n410), .A3(n415), .A4(n420), .Z(data_o[20]) );
  AOI22D0 U499 ( .A1(\data_i[17][21] ), .A2(n683), .B1(\data_i[16][21] ), .B2(
        n684), .ZN(n421) );
  AOI22D0 U500 ( .A1(\data_i[19][21] ), .A2(n685), .B1(\data_i[18][21] ), .B2(
        n686), .ZN(n422) );
  AOI22D0 U501 ( .A1(\data_i[21][21] ), .A2(n687), .B1(\data_i[20][21] ), .B2(
        n688), .ZN(n423) );
  AOI22D0 U502 ( .A1(\data_i[23][21] ), .A2(n689), .B1(\data_i[22][21] ), .B2(
        n690), .ZN(n424) );
  ND4D0 U503 ( .A1(n421), .A2(n422), .A3(n423), .A4(n424), .ZN(n425) );
  AOI22D0 U504 ( .A1(\data_i[25][21] ), .A2(n691), .B1(\data_i[24][21] ), .B2(
        n692), .ZN(n426) );
  AOI22D0 U505 ( .A1(\data_i[27][21] ), .A2(n693), .B1(\data_i[26][21] ), .B2(
        n694), .ZN(n427) );
  AOI22D0 U506 ( .A1(\data_i[29][21] ), .A2(n695), .B1(\data_i[28][21] ), .B2(
        n696), .ZN(n428) );
  AOI22D0 U507 ( .A1(\data_i[31][21] ), .A2(n697), .B1(\data_i[30][21] ), .B2(
        n698), .ZN(n429) );
  ND4D0 U508 ( .A1(n426), .A2(n427), .A3(n428), .A4(n429), .ZN(n430) );
  AOI22D0 U509 ( .A1(\data_i[1][21] ), .A2(n667), .B1(\data_i[0][21] ), .B2(
        n668), .ZN(n431) );
  AOI22D0 U510 ( .A1(\data_i[3][21] ), .A2(n669), .B1(\data_i[2][21] ), .B2(
        n670), .ZN(n432) );
  AOI22D0 U511 ( .A1(\data_i[5][21] ), .A2(n671), .B1(\data_i[4][21] ), .B2(
        n672), .ZN(n433) );
  AOI22D0 U512 ( .A1(\data_i[7][21] ), .A2(n673), .B1(\data_i[6][21] ), .B2(
        n674), .ZN(n434) );
  ND4D0 U513 ( .A1(n431), .A2(n432), .A3(n433), .A4(n434), .ZN(n435) );
  AOI22D0 U514 ( .A1(\data_i[9][21] ), .A2(n675), .B1(\data_i[8][21] ), .B2(
        n676), .ZN(n436) );
  AOI22D0 U515 ( .A1(\data_i[11][21] ), .A2(n677), .B1(\data_i[10][21] ), .B2(
        n678), .ZN(n437) );
  AOI22D0 U516 ( .A1(\data_i[13][21] ), .A2(n679), .B1(\data_i[12][21] ), .B2(
        n680), .ZN(n438) );
  AOI22D0 U517 ( .A1(\data_i[15][21] ), .A2(n681), .B1(\data_i[14][21] ), .B2(
        n682), .ZN(n439) );
  ND4D0 U518 ( .A1(n436), .A2(n437), .A3(n438), .A4(n439), .ZN(n440) );
  OR4D0 U519 ( .A1(n425), .A2(n430), .A3(n435), .A4(n440), .Z(data_o[21]) );
  AOI22D0 U520 ( .A1(\data_i[17][22] ), .A2(n683), .B1(\data_i[16][22] ), .B2(
        n684), .ZN(n441) );
  AOI22D0 U521 ( .A1(\data_i[19][22] ), .A2(n685), .B1(\data_i[18][22] ), .B2(
        n686), .ZN(n442) );
  AOI22D0 U522 ( .A1(\data_i[21][22] ), .A2(n687), .B1(\data_i[20][22] ), .B2(
        n688), .ZN(n443) );
  AOI22D0 U523 ( .A1(\data_i[23][22] ), .A2(n689), .B1(\data_i[22][22] ), .B2(
        n690), .ZN(n444) );
  ND4D0 U524 ( .A1(n441), .A2(n442), .A3(n443), .A4(n444), .ZN(n445) );
  AOI22D0 U525 ( .A1(\data_i[25][22] ), .A2(n691), .B1(\data_i[24][22] ), .B2(
        n692), .ZN(n446) );
  AOI22D0 U526 ( .A1(\data_i[27][22] ), .A2(n693), .B1(\data_i[26][22] ), .B2(
        n694), .ZN(n447) );
  AOI22D0 U527 ( .A1(\data_i[29][22] ), .A2(n695), .B1(\data_i[28][22] ), .B2(
        n696), .ZN(n448) );
  AOI22D0 U528 ( .A1(\data_i[31][22] ), .A2(n697), .B1(\data_i[30][22] ), .B2(
        n698), .ZN(n449) );
  ND4D0 U529 ( .A1(n446), .A2(n447), .A3(n448), .A4(n449), .ZN(n450) );
  AOI22D0 U530 ( .A1(\data_i[1][22] ), .A2(n667), .B1(\data_i[0][22] ), .B2(
        n668), .ZN(n451) );
  AOI22D0 U531 ( .A1(\data_i[3][22] ), .A2(n669), .B1(\data_i[2][22] ), .B2(
        n670), .ZN(n452) );
  AOI22D0 U532 ( .A1(\data_i[5][22] ), .A2(n671), .B1(\data_i[4][22] ), .B2(
        n672), .ZN(n453) );
  AOI22D0 U533 ( .A1(\data_i[7][22] ), .A2(n673), .B1(\data_i[6][22] ), .B2(
        n674), .ZN(n454) );
  ND4D0 U534 ( .A1(n451), .A2(n452), .A3(n453), .A4(n454), .ZN(n455) );
  AOI22D0 U535 ( .A1(\data_i[9][22] ), .A2(n675), .B1(\data_i[8][22] ), .B2(
        n676), .ZN(n456) );
  AOI22D0 U536 ( .A1(\data_i[11][22] ), .A2(n677), .B1(\data_i[10][22] ), .B2(
        n678), .ZN(n457) );
  AOI22D0 U537 ( .A1(\data_i[13][22] ), .A2(n679), .B1(\data_i[12][22] ), .B2(
        n680), .ZN(n458) );
  AOI22D0 U538 ( .A1(\data_i[15][22] ), .A2(n681), .B1(\data_i[14][22] ), .B2(
        n682), .ZN(n459) );
  ND4D0 U539 ( .A1(n456), .A2(n457), .A3(n458), .A4(n459), .ZN(n460) );
  OR4D0 U540 ( .A1(n445), .A2(n450), .A3(n455), .A4(n460), .Z(data_o[22]) );
  AOI22D0 U541 ( .A1(\data_i[17][23] ), .A2(n683), .B1(\data_i[16][23] ), .B2(
        n684), .ZN(n461) );
  AOI22D0 U542 ( .A1(\data_i[19][23] ), .A2(n685), .B1(\data_i[18][23] ), .B2(
        n686), .ZN(n462) );
  AOI22D0 U543 ( .A1(\data_i[21][23] ), .A2(n687), .B1(\data_i[20][23] ), .B2(
        n688), .ZN(n463) );
  AOI22D0 U544 ( .A1(\data_i[23][23] ), .A2(n689), .B1(\data_i[22][23] ), .B2(
        n690), .ZN(n464) );
  ND4D0 U545 ( .A1(n461), .A2(n462), .A3(n463), .A4(n464), .ZN(n465) );
  AOI22D0 U546 ( .A1(\data_i[25][23] ), .A2(n691), .B1(\data_i[24][23] ), .B2(
        n692), .ZN(n466) );
  AOI22D0 U547 ( .A1(\data_i[27][23] ), .A2(n693), .B1(\data_i[26][23] ), .B2(
        n694), .ZN(n467) );
  AOI22D0 U548 ( .A1(\data_i[29][23] ), .A2(n695), .B1(\data_i[28][23] ), .B2(
        n696), .ZN(n468) );
  AOI22D0 U549 ( .A1(\data_i[31][23] ), .A2(n697), .B1(\data_i[30][23] ), .B2(
        n698), .ZN(n469) );
  ND4D0 U550 ( .A1(n466), .A2(n467), .A3(n468), .A4(n469), .ZN(n470) );
  AOI22D0 U551 ( .A1(\data_i[1][23] ), .A2(n667), .B1(\data_i[0][23] ), .B2(
        n668), .ZN(n471) );
  AOI22D0 U552 ( .A1(\data_i[3][23] ), .A2(n669), .B1(\data_i[2][23] ), .B2(
        n670), .ZN(n472) );
  AOI22D0 U553 ( .A1(\data_i[5][23] ), .A2(n671), .B1(\data_i[4][23] ), .B2(
        n672), .ZN(n473) );
  AOI22D0 U554 ( .A1(\data_i[7][23] ), .A2(n673), .B1(\data_i[6][23] ), .B2(
        n674), .ZN(n474) );
  ND4D0 U555 ( .A1(n471), .A2(n472), .A3(n473), .A4(n474), .ZN(n475) );
  AOI22D0 U556 ( .A1(\data_i[9][23] ), .A2(n675), .B1(\data_i[8][23] ), .B2(
        n676), .ZN(n476) );
  AOI22D0 U557 ( .A1(\data_i[11][23] ), .A2(n677), .B1(\data_i[10][23] ), .B2(
        n678), .ZN(n477) );
  AOI22D0 U558 ( .A1(\data_i[13][23] ), .A2(n679), .B1(\data_i[12][23] ), .B2(
        n680), .ZN(n478) );
  AOI22D0 U559 ( .A1(\data_i[15][23] ), .A2(n681), .B1(\data_i[14][23] ), .B2(
        n682), .ZN(n479) );
  ND4D0 U560 ( .A1(n476), .A2(n477), .A3(n478), .A4(n479), .ZN(n480) );
  OR4D0 U561 ( .A1(n465), .A2(n470), .A3(n475), .A4(n480), .Z(data_o[23]) );
  AOI22D0 U562 ( .A1(\data_i[17][24] ), .A2(n683), .B1(\data_i[16][24] ), .B2(
        n684), .ZN(n481) );
  AOI22D0 U563 ( .A1(\data_i[19][24] ), .A2(n685), .B1(\data_i[18][24] ), .B2(
        n686), .ZN(n482) );
  AOI22D0 U564 ( .A1(\data_i[21][24] ), .A2(n687), .B1(\data_i[20][24] ), .B2(
        n688), .ZN(n483) );
  AOI22D0 U565 ( .A1(\data_i[23][24] ), .A2(n689), .B1(\data_i[22][24] ), .B2(
        n690), .ZN(n484) );
  ND4D0 U566 ( .A1(n481), .A2(n482), .A3(n483), .A4(n484), .ZN(n485) );
  AOI22D0 U567 ( .A1(\data_i[25][24] ), .A2(n691), .B1(\data_i[24][24] ), .B2(
        n692), .ZN(n486) );
  AOI22D0 U568 ( .A1(\data_i[27][24] ), .A2(n693), .B1(\data_i[26][24] ), .B2(
        n694), .ZN(n487) );
  AOI22D0 U569 ( .A1(\data_i[29][24] ), .A2(n695), .B1(\data_i[28][24] ), .B2(
        n696), .ZN(n488) );
  AOI22D0 U570 ( .A1(\data_i[31][24] ), .A2(n697), .B1(\data_i[30][24] ), .B2(
        n698), .ZN(n489) );
  ND4D0 U571 ( .A1(n486), .A2(n487), .A3(n488), .A4(n489), .ZN(n490) );
  AOI22D0 U572 ( .A1(\data_i[1][24] ), .A2(n667), .B1(\data_i[0][24] ), .B2(
        n668), .ZN(n491) );
  AOI22D0 U573 ( .A1(\data_i[3][24] ), .A2(n669), .B1(\data_i[2][24] ), .B2(
        n670), .ZN(n492) );
  AOI22D0 U574 ( .A1(\data_i[5][24] ), .A2(n671), .B1(\data_i[4][24] ), .B2(
        n672), .ZN(n493) );
  AOI22D0 U575 ( .A1(\data_i[7][24] ), .A2(n673), .B1(\data_i[6][24] ), .B2(
        n674), .ZN(n494) );
  ND4D0 U576 ( .A1(n491), .A2(n492), .A3(n493), .A4(n494), .ZN(n495) );
  AOI22D0 U577 ( .A1(\data_i[9][24] ), .A2(n675), .B1(\data_i[8][24] ), .B2(
        n676), .ZN(n496) );
  AOI22D0 U578 ( .A1(\data_i[11][24] ), .A2(n677), .B1(\data_i[10][24] ), .B2(
        n678), .ZN(n497) );
  AOI22D0 U579 ( .A1(\data_i[13][24] ), .A2(n679), .B1(\data_i[12][24] ), .B2(
        n680), .ZN(n498) );
  AOI22D0 U580 ( .A1(\data_i[15][24] ), .A2(n681), .B1(\data_i[14][24] ), .B2(
        n682), .ZN(n499) );
  ND4D0 U581 ( .A1(n496), .A2(n497), .A3(n498), .A4(n499), .ZN(n500) );
  OR4D0 U582 ( .A1(n485), .A2(n490), .A3(n495), .A4(n500), .Z(data_o[24]) );
  AOI22D0 U583 ( .A1(\data_i[17][25] ), .A2(n683), .B1(\data_i[16][25] ), .B2(
        n684), .ZN(n501) );
  AOI22D0 U584 ( .A1(\data_i[19][25] ), .A2(n685), .B1(\data_i[18][25] ), .B2(
        n686), .ZN(n502) );
  AOI22D0 U585 ( .A1(\data_i[21][25] ), .A2(n687), .B1(\data_i[20][25] ), .B2(
        n688), .ZN(n503) );
  AOI22D0 U586 ( .A1(\data_i[23][25] ), .A2(n689), .B1(\data_i[22][25] ), .B2(
        n690), .ZN(n504) );
  ND4D0 U587 ( .A1(n501), .A2(n502), .A3(n503), .A4(n504), .ZN(n505) );
  AOI22D0 U588 ( .A1(\data_i[25][25] ), .A2(n691), .B1(\data_i[24][25] ), .B2(
        n692), .ZN(n506) );
  AOI22D0 U589 ( .A1(\data_i[27][25] ), .A2(n693), .B1(\data_i[26][25] ), .B2(
        n694), .ZN(n507) );
  AOI22D0 U590 ( .A1(\data_i[29][25] ), .A2(n695), .B1(\data_i[28][25] ), .B2(
        n696), .ZN(n508) );
  AOI22D0 U591 ( .A1(\data_i[31][25] ), .A2(n697), .B1(\data_i[30][25] ), .B2(
        n698), .ZN(n509) );
  ND4D0 U592 ( .A1(n506), .A2(n507), .A3(n508), .A4(n509), .ZN(n510) );
  AOI22D0 U593 ( .A1(\data_i[1][25] ), .A2(n667), .B1(\data_i[0][25] ), .B2(
        n668), .ZN(n511) );
  AOI22D0 U594 ( .A1(\data_i[3][25] ), .A2(n669), .B1(\data_i[2][25] ), .B2(
        n670), .ZN(n512) );
  AOI22D0 U595 ( .A1(\data_i[5][25] ), .A2(n671), .B1(\data_i[4][25] ), .B2(
        n672), .ZN(n513) );
  AOI22D0 U596 ( .A1(\data_i[7][25] ), .A2(n673), .B1(\data_i[6][25] ), .B2(
        n674), .ZN(n514) );
  ND4D0 U597 ( .A1(n511), .A2(n512), .A3(n513), .A4(n514), .ZN(n515) );
  AOI22D0 U598 ( .A1(\data_i[9][25] ), .A2(n675), .B1(\data_i[8][25] ), .B2(
        n676), .ZN(n516) );
  AOI22D0 U599 ( .A1(\data_i[11][25] ), .A2(n677), .B1(\data_i[10][25] ), .B2(
        n678), .ZN(n517) );
  AOI22D0 U600 ( .A1(\data_i[13][25] ), .A2(n679), .B1(\data_i[12][25] ), .B2(
        n680), .ZN(n518) );
  AOI22D0 U601 ( .A1(\data_i[15][25] ), .A2(n681), .B1(\data_i[14][25] ), .B2(
        n682), .ZN(n519) );
  ND4D0 U602 ( .A1(n516), .A2(n517), .A3(n518), .A4(n519), .ZN(n520) );
  OR4D0 U603 ( .A1(n505), .A2(n510), .A3(n515), .A4(n520), .Z(data_o[25]) );
  AOI22D0 U604 ( .A1(\data_i[17][26] ), .A2(n683), .B1(\data_i[16][26] ), .B2(
        n684), .ZN(n521) );
  AOI22D0 U605 ( .A1(\data_i[19][26] ), .A2(n685), .B1(\data_i[18][26] ), .B2(
        n686), .ZN(n522) );
  AOI22D0 U606 ( .A1(\data_i[21][26] ), .A2(n687), .B1(\data_i[20][26] ), .B2(
        n688), .ZN(n523) );
  AOI22D0 U607 ( .A1(\data_i[23][26] ), .A2(n689), .B1(\data_i[22][26] ), .B2(
        n690), .ZN(n524) );
  ND4D0 U608 ( .A1(n521), .A2(n522), .A3(n523), .A4(n524), .ZN(n525) );
  AOI22D0 U609 ( .A1(\data_i[25][26] ), .A2(n691), .B1(\data_i[24][26] ), .B2(
        n692), .ZN(n526) );
  AOI22D0 U610 ( .A1(\data_i[27][26] ), .A2(n693), .B1(\data_i[26][26] ), .B2(
        n694), .ZN(n527) );
  AOI22D0 U611 ( .A1(\data_i[29][26] ), .A2(n695), .B1(\data_i[28][26] ), .B2(
        n696), .ZN(n528) );
  AOI22D0 U612 ( .A1(\data_i[31][26] ), .A2(n697), .B1(\data_i[30][26] ), .B2(
        n698), .ZN(n529) );
  ND4D0 U613 ( .A1(n526), .A2(n527), .A3(n528), .A4(n529), .ZN(n530) );
  AOI22D0 U614 ( .A1(\data_i[1][26] ), .A2(n667), .B1(\data_i[0][26] ), .B2(
        n668), .ZN(n531) );
  AOI22D0 U615 ( .A1(\data_i[3][26] ), .A2(n669), .B1(\data_i[2][26] ), .B2(
        n670), .ZN(n532) );
  AOI22D0 U616 ( .A1(\data_i[5][26] ), .A2(n671), .B1(\data_i[4][26] ), .B2(
        n672), .ZN(n533) );
  AOI22D0 U617 ( .A1(\data_i[7][26] ), .A2(n673), .B1(\data_i[6][26] ), .B2(
        n674), .ZN(n534) );
  ND4D0 U618 ( .A1(n531), .A2(n532), .A3(n533), .A4(n534), .ZN(n535) );
  AOI22D0 U619 ( .A1(\data_i[9][26] ), .A2(n675), .B1(\data_i[8][26] ), .B2(
        n676), .ZN(n536) );
  AOI22D0 U620 ( .A1(\data_i[11][26] ), .A2(n677), .B1(\data_i[10][26] ), .B2(
        n678), .ZN(n537) );
  AOI22D0 U621 ( .A1(\data_i[13][26] ), .A2(n679), .B1(\data_i[12][26] ), .B2(
        n680), .ZN(n538) );
  AOI22D0 U622 ( .A1(\data_i[15][26] ), .A2(n681), .B1(\data_i[14][26] ), .B2(
        n682), .ZN(n539) );
  ND4D0 U623 ( .A1(n536), .A2(n537), .A3(n538), .A4(n539), .ZN(n540) );
  OR4D0 U624 ( .A1(n525), .A2(n530), .A3(n535), .A4(n540), .Z(data_o[26]) );
  AOI22D0 U625 ( .A1(\data_i[17][27] ), .A2(n683), .B1(\data_i[16][27] ), .B2(
        n684), .ZN(n541) );
  AOI22D0 U626 ( .A1(\data_i[19][27] ), .A2(n685), .B1(\data_i[18][27] ), .B2(
        n686), .ZN(n542) );
  AOI22D0 U627 ( .A1(\data_i[21][27] ), .A2(n687), .B1(\data_i[20][27] ), .B2(
        n688), .ZN(n543) );
  AOI22D0 U628 ( .A1(\data_i[23][27] ), .A2(n689), .B1(\data_i[22][27] ), .B2(
        n690), .ZN(n544) );
  ND4D0 U629 ( .A1(n541), .A2(n542), .A3(n543), .A4(n544), .ZN(n545) );
  AOI22D0 U630 ( .A1(\data_i[25][27] ), .A2(n691), .B1(\data_i[24][27] ), .B2(
        n692), .ZN(n546) );
  AOI22D0 U631 ( .A1(\data_i[27][27] ), .A2(n693), .B1(\data_i[26][27] ), .B2(
        n694), .ZN(n547) );
  AOI22D0 U632 ( .A1(\data_i[29][27] ), .A2(n695), .B1(\data_i[28][27] ), .B2(
        n696), .ZN(n548) );
  AOI22D0 U633 ( .A1(\data_i[31][27] ), .A2(n697), .B1(\data_i[30][27] ), .B2(
        n698), .ZN(n549) );
  ND4D0 U634 ( .A1(n546), .A2(n547), .A3(n548), .A4(n549), .ZN(n550) );
  AOI22D0 U635 ( .A1(\data_i[1][27] ), .A2(n667), .B1(\data_i[0][27] ), .B2(
        n668), .ZN(n551) );
  AOI22D0 U636 ( .A1(\data_i[3][27] ), .A2(n669), .B1(\data_i[2][27] ), .B2(
        n670), .ZN(n552) );
  AOI22D0 U637 ( .A1(\data_i[5][27] ), .A2(n671), .B1(\data_i[4][27] ), .B2(
        n672), .ZN(n553) );
  AOI22D0 U638 ( .A1(\data_i[7][27] ), .A2(n673), .B1(\data_i[6][27] ), .B2(
        n674), .ZN(n554) );
  ND4D0 U639 ( .A1(n551), .A2(n552), .A3(n553), .A4(n554), .ZN(n555) );
  AOI22D0 U640 ( .A1(\data_i[9][27] ), .A2(n675), .B1(\data_i[8][27] ), .B2(
        n676), .ZN(n556) );
  AOI22D0 U641 ( .A1(\data_i[11][27] ), .A2(n677), .B1(\data_i[10][27] ), .B2(
        n678), .ZN(n557) );
  AOI22D0 U642 ( .A1(\data_i[13][27] ), .A2(n679), .B1(\data_i[12][27] ), .B2(
        n680), .ZN(n558) );
  AOI22D0 U643 ( .A1(\data_i[15][27] ), .A2(n681), .B1(\data_i[14][27] ), .B2(
        n682), .ZN(n559) );
  ND4D0 U644 ( .A1(n556), .A2(n557), .A3(n558), .A4(n559), .ZN(n560) );
  OR4D0 U645 ( .A1(n545), .A2(n550), .A3(n555), .A4(n560), .Z(data_o[27]) );
  AOI22D0 U646 ( .A1(\data_i[17][28] ), .A2(n683), .B1(\data_i[16][28] ), .B2(
        n684), .ZN(n561) );
  AOI22D0 U647 ( .A1(\data_i[19][28] ), .A2(n685), .B1(\data_i[18][28] ), .B2(
        n686), .ZN(n562) );
  AOI22D0 U648 ( .A1(\data_i[21][28] ), .A2(n687), .B1(\data_i[20][28] ), .B2(
        n688), .ZN(n563) );
  AOI22D0 U649 ( .A1(\data_i[23][28] ), .A2(n689), .B1(\data_i[22][28] ), .B2(
        n690), .ZN(n564) );
  ND4D0 U650 ( .A1(n561), .A2(n562), .A3(n563), .A4(n564), .ZN(n565) );
  AOI22D0 U651 ( .A1(\data_i[25][28] ), .A2(n691), .B1(\data_i[24][28] ), .B2(
        n692), .ZN(n566) );
  AOI22D0 U652 ( .A1(\data_i[27][28] ), .A2(n693), .B1(\data_i[26][28] ), .B2(
        n694), .ZN(n567) );
  AOI22D0 U653 ( .A1(\data_i[29][28] ), .A2(n695), .B1(\data_i[28][28] ), .B2(
        n696), .ZN(n568) );
  AOI22D0 U654 ( .A1(\data_i[31][28] ), .A2(n697), .B1(\data_i[30][28] ), .B2(
        n698), .ZN(n569) );
  ND4D0 U655 ( .A1(n566), .A2(n567), .A3(n568), .A4(n569), .ZN(n570) );
  AOI22D0 U656 ( .A1(\data_i[1][28] ), .A2(n667), .B1(\data_i[0][28] ), .B2(
        n668), .ZN(n571) );
  AOI22D0 U657 ( .A1(\data_i[3][28] ), .A2(n669), .B1(\data_i[2][28] ), .B2(
        n670), .ZN(n572) );
  AOI22D0 U658 ( .A1(\data_i[5][28] ), .A2(n671), .B1(\data_i[4][28] ), .B2(
        n672), .ZN(n573) );
  AOI22D0 U659 ( .A1(\data_i[7][28] ), .A2(n673), .B1(\data_i[6][28] ), .B2(
        n674), .ZN(n574) );
  ND4D0 U660 ( .A1(n571), .A2(n572), .A3(n573), .A4(n574), .ZN(n575) );
  AOI22D0 U661 ( .A1(\data_i[9][28] ), .A2(n675), .B1(\data_i[8][28] ), .B2(
        n676), .ZN(n576) );
  AOI22D0 U662 ( .A1(\data_i[11][28] ), .A2(n677), .B1(\data_i[10][28] ), .B2(
        n678), .ZN(n577) );
  AOI22D0 U663 ( .A1(\data_i[13][28] ), .A2(n679), .B1(\data_i[12][28] ), .B2(
        n680), .ZN(n578) );
  AOI22D0 U664 ( .A1(\data_i[15][28] ), .A2(n681), .B1(\data_i[14][28] ), .B2(
        n682), .ZN(n579) );
  ND4D0 U665 ( .A1(n576), .A2(n577), .A3(n578), .A4(n579), .ZN(n580) );
  OR4D0 U666 ( .A1(n565), .A2(n570), .A3(n575), .A4(n580), .Z(data_o[28]) );
  AOI22D0 U667 ( .A1(\data_i[17][29] ), .A2(n683), .B1(\data_i[16][29] ), .B2(
        n684), .ZN(n581) );
  AOI22D0 U668 ( .A1(\data_i[19][29] ), .A2(n685), .B1(\data_i[18][29] ), .B2(
        n686), .ZN(n582) );
  AOI22D0 U669 ( .A1(\data_i[21][29] ), .A2(n687), .B1(\data_i[20][29] ), .B2(
        n688), .ZN(n583) );
  AOI22D0 U670 ( .A1(\data_i[23][29] ), .A2(n689), .B1(\data_i[22][29] ), .B2(
        n690), .ZN(n584) );
  ND4D0 U671 ( .A1(n581), .A2(n582), .A3(n583), .A4(n584), .ZN(n585) );
  AOI22D0 U672 ( .A1(\data_i[25][29] ), .A2(n691), .B1(\data_i[24][29] ), .B2(
        n692), .ZN(n586) );
  AOI22D0 U673 ( .A1(\data_i[27][29] ), .A2(n693), .B1(\data_i[26][29] ), .B2(
        n694), .ZN(n587) );
  AOI22D0 U674 ( .A1(\data_i[29][29] ), .A2(n695), .B1(\data_i[28][29] ), .B2(
        n696), .ZN(n588) );
  AOI22D0 U675 ( .A1(\data_i[31][29] ), .A2(n697), .B1(\data_i[30][29] ), .B2(
        n698), .ZN(n589) );
  ND4D0 U676 ( .A1(n586), .A2(n587), .A3(n588), .A4(n589), .ZN(n590) );
  AOI22D0 U677 ( .A1(\data_i[1][29] ), .A2(n667), .B1(\data_i[0][29] ), .B2(
        n668), .ZN(n591) );
  AOI22D0 U678 ( .A1(\data_i[3][29] ), .A2(n669), .B1(\data_i[2][29] ), .B2(
        n670), .ZN(n592) );
  AOI22D0 U679 ( .A1(\data_i[5][29] ), .A2(n671), .B1(\data_i[4][29] ), .B2(
        n672), .ZN(n593) );
  AOI22D0 U680 ( .A1(\data_i[7][29] ), .A2(n673), .B1(\data_i[6][29] ), .B2(
        n674), .ZN(n594) );
  ND4D0 U681 ( .A1(n591), .A2(n592), .A3(n593), .A4(n594), .ZN(n595) );
  AOI22D0 U682 ( .A1(\data_i[9][29] ), .A2(n675), .B1(\data_i[8][29] ), .B2(
        n676), .ZN(n596) );
  AOI22D0 U683 ( .A1(\data_i[11][29] ), .A2(n677), .B1(\data_i[10][29] ), .B2(
        n678), .ZN(n597) );
  AOI22D0 U684 ( .A1(\data_i[13][29] ), .A2(n679), .B1(\data_i[12][29] ), .B2(
        n680), .ZN(n598) );
  AOI22D0 U685 ( .A1(\data_i[15][29] ), .A2(n681), .B1(\data_i[14][29] ), .B2(
        n682), .ZN(n599) );
  ND4D0 U686 ( .A1(n596), .A2(n597), .A3(n598), .A4(n599), .ZN(n600) );
  OR4D0 U687 ( .A1(n585), .A2(n590), .A3(n595), .A4(n600), .Z(data_o[29]) );
  AOI22D0 U688 ( .A1(\data_i[17][30] ), .A2(n683), .B1(\data_i[16][30] ), .B2(
        n684), .ZN(n601) );
  AOI22D0 U689 ( .A1(\data_i[19][30] ), .A2(n685), .B1(\data_i[18][30] ), .B2(
        n686), .ZN(n602) );
  AOI22D0 U690 ( .A1(\data_i[21][30] ), .A2(n687), .B1(\data_i[20][30] ), .B2(
        n688), .ZN(n603) );
  AOI22D0 U691 ( .A1(\data_i[23][30] ), .A2(n689), .B1(\data_i[22][30] ), .B2(
        n690), .ZN(n604) );
  ND4D0 U692 ( .A1(n601), .A2(n602), .A3(n603), .A4(n604), .ZN(n605) );
  AOI22D0 U693 ( .A1(\data_i[25][30] ), .A2(n691), .B1(\data_i[24][30] ), .B2(
        n692), .ZN(n606) );
  AOI22D0 U694 ( .A1(\data_i[27][30] ), .A2(n693), .B1(\data_i[26][30] ), .B2(
        n694), .ZN(n607) );
  AOI22D0 U695 ( .A1(\data_i[29][30] ), .A2(n695), .B1(\data_i[28][30] ), .B2(
        n696), .ZN(n608) );
  AOI22D0 U696 ( .A1(\data_i[31][30] ), .A2(n697), .B1(\data_i[30][30] ), .B2(
        n698), .ZN(n609) );
  ND4D0 U697 ( .A1(n606), .A2(n607), .A3(n608), .A4(n609), .ZN(n610) );
  AOI22D0 U698 ( .A1(\data_i[1][30] ), .A2(n667), .B1(\data_i[0][30] ), .B2(
        n668), .ZN(n611) );
  AOI22D0 U699 ( .A1(\data_i[3][30] ), .A2(n669), .B1(\data_i[2][30] ), .B2(
        n670), .ZN(n612) );
  AOI22D0 U700 ( .A1(\data_i[5][30] ), .A2(n671), .B1(\data_i[4][30] ), .B2(
        n672), .ZN(n613) );
  AOI22D0 U701 ( .A1(\data_i[7][30] ), .A2(n673), .B1(\data_i[6][30] ), .B2(
        n674), .ZN(n614) );
  ND4D0 U702 ( .A1(n611), .A2(n612), .A3(n613), .A4(n614), .ZN(n615) );
  AOI22D0 U703 ( .A1(\data_i[9][30] ), .A2(n675), .B1(\data_i[8][30] ), .B2(
        n676), .ZN(n616) );
  AOI22D0 U704 ( .A1(\data_i[11][30] ), .A2(n677), .B1(\data_i[10][30] ), .B2(
        n678), .ZN(n617) );
  AOI22D0 U705 ( .A1(\data_i[13][30] ), .A2(n679), .B1(\data_i[12][30] ), .B2(
        n680), .ZN(n618) );
  AOI22D0 U706 ( .A1(\data_i[15][30] ), .A2(n681), .B1(\data_i[14][30] ), .B2(
        n682), .ZN(n619) );
  ND4D0 U707 ( .A1(n616), .A2(n617), .A3(n618), .A4(n619), .ZN(n620) );
  OR4D0 U708 ( .A1(n605), .A2(n610), .A3(n615), .A4(n620), .Z(data_o[30]) );
  AOI22D0 U709 ( .A1(\data_i[17][31] ), .A2(n683), .B1(\data_i[16][31] ), .B2(
        n684), .ZN(n621) );
  AOI22D0 U710 ( .A1(\data_i[19][31] ), .A2(n685), .B1(\data_i[18][31] ), .B2(
        n686), .ZN(n622) );
  AOI22D0 U711 ( .A1(\data_i[21][31] ), .A2(n687), .B1(\data_i[20][31] ), .B2(
        n688), .ZN(n623) );
  AOI22D0 U712 ( .A1(\data_i[23][31] ), .A2(n689), .B1(\data_i[22][31] ), .B2(
        n690), .ZN(n624) );
  ND4D0 U713 ( .A1(n621), .A2(n622), .A3(n623), .A4(n624), .ZN(n625) );
  AOI22D0 U714 ( .A1(\data_i[25][31] ), .A2(n691), .B1(\data_i[24][31] ), .B2(
        n692), .ZN(n626) );
  AOI22D0 U715 ( .A1(\data_i[27][31] ), .A2(n693), .B1(\data_i[26][31] ), .B2(
        n694), .ZN(n627) );
  AOI22D0 U716 ( .A1(\data_i[29][31] ), .A2(n695), .B1(\data_i[28][31] ), .B2(
        n696), .ZN(n628) );
  AOI22D0 U717 ( .A1(\data_i[31][31] ), .A2(n697), .B1(\data_i[30][31] ), .B2(
        n698), .ZN(n629) );
  ND4D0 U718 ( .A1(n626), .A2(n627), .A3(n628), .A4(n629), .ZN(n630) );
  AOI22D0 U719 ( .A1(\data_i[1][31] ), .A2(n667), .B1(\data_i[0][31] ), .B2(
        n668), .ZN(n631) );
  AOI22D0 U720 ( .A1(\data_i[3][31] ), .A2(n669), .B1(\data_i[2][31] ), .B2(
        n670), .ZN(n632) );
  AOI22D0 U721 ( .A1(\data_i[5][31] ), .A2(n671), .B1(\data_i[4][31] ), .B2(
        n672), .ZN(n633) );
  AOI22D0 U722 ( .A1(\data_i[7][31] ), .A2(n673), .B1(\data_i[6][31] ), .B2(
        n674), .ZN(n634) );
  ND4D0 U723 ( .A1(n631), .A2(n632), .A3(n633), .A4(n634), .ZN(n635) );
  AOI22D0 U724 ( .A1(\data_i[9][31] ), .A2(n675), .B1(\data_i[8][31] ), .B2(
        n676), .ZN(n636) );
  AOI22D0 U725 ( .A1(\data_i[11][31] ), .A2(n677), .B1(\data_i[10][31] ), .B2(
        n678), .ZN(n637) );
  AOI22D0 U726 ( .A1(\data_i[13][31] ), .A2(n679), .B1(\data_i[12][31] ), .B2(
        n680), .ZN(n638) );
  AOI22D0 U727 ( .A1(\data_i[15][31] ), .A2(n681), .B1(\data_i[14][31] ), .B2(
        n682), .ZN(n639) );
  ND4D0 U728 ( .A1(n636), .A2(n637), .A3(n638), .A4(n639), .ZN(n640) );
  OR4D0 U729 ( .A1(n625), .A2(n630), .A3(n635), .A4(n640), .Z(data_o[31]) );
  ND2D1 U730 ( .A1(select_i[4]), .A2(n652), .ZN(n659) );
endmodule


module decoder_5_32_0 ( decoder_i, decoder_o );
  input [4:0] decoder_i;
  output [31:0] decoder_o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;

  NR2D1 U1 ( .A1(decoder_i[0]), .A2(n8), .ZN(n7) );
  INVD1 U2 ( .I(decoder_i[1]), .ZN(n8) );
  INVD1 U3 ( .I(decoder_i[4]), .ZN(n9) );
  NR2D1 U4 ( .A1(decoder_i[1]), .A2(decoder_i[0]), .ZN(n10) );
  INVD1 U5 ( .I(decoder_i[2]), .ZN(n1) );
  INVD1 U6 ( .I(decoder_i[3]), .ZN(n2) );
  ND3D1 U7 ( .A1(decoder_i[4]), .A2(decoder_i[1]), .A3(decoder_i[0]), .ZN(n3)
         );
  ND2D1 U8 ( .A1(decoder_i[4]), .A2(n7), .ZN(n4) );
  ND3D1 U9 ( .A1(decoder_i[4]), .A2(decoder_i[0]), .A3(n8), .ZN(n5) );
  ND2D1 U10 ( .A1(decoder_i[4]), .A2(n10), .ZN(n6) );
  ND2D1 U11 ( .A1(decoder_i[3]), .A2(decoder_i[2]), .ZN(n11) );
  ND2D1 U12 ( .A1(decoder_i[3]), .A2(n1), .ZN(n12) );
  ND2D1 U13 ( .A1(decoder_i[2]), .A2(n2), .ZN(n13) );
  ND3D1 U14 ( .A1(decoder_i[1]), .A2(decoder_i[0]), .A3(n9), .ZN(n14) );
  ND2D1 U15 ( .A1(n7), .A2(n9), .ZN(n15) );
  ND3D1 U16 ( .A1(decoder_i[0]), .A2(n9), .A3(n8), .ZN(n16) );
  ND2D1 U17 ( .A1(n10), .A2(n9), .ZN(n17) );
  ND2D1 U18 ( .A1(n2), .A2(n1), .ZN(n18) );
  NR2D1 U19 ( .A1(n11), .A2(n3), .ZN(decoder_o[31]) );
  NR2D1 U20 ( .A1(n11), .A2(n6), .ZN(decoder_o[28]) );
  NR2D1 U21 ( .A1(n11), .A2(n17), .ZN(decoder_o[12]) );
  NR2D1 U22 ( .A1(n12), .A2(n17), .ZN(decoder_o[8]) );
  NR2D1 U23 ( .A1(n18), .A2(n17), .ZN(decoder_o[0]) );
  NR2D1 U24 ( .A1(n6), .A2(n12), .ZN(decoder_o[24]) );
  NR2D1 U25 ( .A1(n6), .A2(n18), .ZN(decoder_o[16]) );
  NR2D1 U26 ( .A1(n13), .A2(n17), .ZN(decoder_o[4]) );
  NR2D1 U27 ( .A1(n6), .A2(n13), .ZN(decoder_o[20]) );
  NR2D1 U28 ( .A1(n3), .A2(n12), .ZN(decoder_o[27]) );
  NR2D1 U29 ( .A1(n3), .A2(n18), .ZN(decoder_o[19]) );
  NR2D1 U30 ( .A1(n3), .A2(n13), .ZN(decoder_o[23]) );
  NR2D1 U31 ( .A1(n5), .A2(n13), .ZN(decoder_o[21]) );
  NR2D1 U32 ( .A1(n5), .A2(n12), .ZN(decoder_o[25]) );
  NR2D1 U33 ( .A1(n5), .A2(n18), .ZN(decoder_o[17]) );
  NR2D1 U34 ( .A1(n11), .A2(n5), .ZN(decoder_o[29]) );
  NR2D1 U35 ( .A1(n11), .A2(n16), .ZN(decoder_o[13]) );
  NR2D1 U36 ( .A1(n18), .A2(n16), .ZN(decoder_o[1]) );
  NR2D1 U37 ( .A1(n13), .A2(n16), .ZN(decoder_o[5]) );
  NR2D1 U38 ( .A1(n12), .A2(n16), .ZN(decoder_o[9]) );
  NR2D1 U39 ( .A1(n11), .A2(n14), .ZN(decoder_o[15]) );
  NR2D1 U40 ( .A1(n18), .A2(n14), .ZN(decoder_o[3]) );
  NR2D1 U41 ( .A1(n12), .A2(n14), .ZN(decoder_o[11]) );
  NR2D1 U42 ( .A1(n13), .A2(n14), .ZN(decoder_o[7]) );
  NR2D1 U43 ( .A1(n4), .A2(n12), .ZN(decoder_o[26]) );
  NR2D1 U44 ( .A1(n4), .A2(n18), .ZN(decoder_o[18]) );
  NR2D1 U45 ( .A1(n4), .A2(n13), .ZN(decoder_o[22]) );
  NR2D1 U46 ( .A1(n11), .A2(n4), .ZN(decoder_o[30]) );
  NR2D1 U47 ( .A1(n11), .A2(n15), .ZN(decoder_o[14]) );
  NR2D1 U48 ( .A1(n12), .A2(n15), .ZN(decoder_o[10]) );
  NR2D1 U49 ( .A1(n13), .A2(n15), .ZN(decoder_o[6]) );
  NR2D1 U50 ( .A1(n18), .A2(n15), .ZN(decoder_o[2]) );
endmodule


module cam ( reset, clk, read, read_index, write, write_index, write_data, 
        search, search_data, read_valid, read_value, search_valid, 
        search_index );
  input [4:0] read_index;
  input [4:0] write_index;
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  output [4:0] search_index;
  input reset, clk, read, write, search;
  output read_valid, search_valid;
  wire   \read_value_mux[31][31] , \read_value_mux[31][30] ,
         \read_value_mux[31][29] , \read_value_mux[31][28] ,
         \read_value_mux[31][27] , \read_value_mux[31][26] ,
         \read_value_mux[31][25] , \read_value_mux[31][24] ,
         \read_value_mux[31][23] , \read_value_mux[31][22] ,
         \read_value_mux[31][21] , \read_value_mux[31][20] ,
         \read_value_mux[31][19] , \read_value_mux[31][18] ,
         \read_value_mux[31][17] , \read_value_mux[31][16] ,
         \read_value_mux[31][15] , \read_value_mux[31][14] ,
         \read_value_mux[31][13] , \read_value_mux[31][12] ,
         \read_value_mux[31][11] , \read_value_mux[31][10] ,
         \read_value_mux[31][9] , \read_value_mux[31][8] ,
         \read_value_mux[31][7] , \read_value_mux[31][6] ,
         \read_value_mux[31][5] , \read_value_mux[31][4] ,
         \read_value_mux[31][3] , \read_value_mux[31][2] ,
         \read_value_mux[31][1] , \read_value_mux[31][0] ,
         \read_value_mux[30][31] , \read_value_mux[30][30] ,
         \read_value_mux[30][29] , \read_value_mux[30][28] ,
         \read_value_mux[30][27] , \read_value_mux[30][26] ,
         \read_value_mux[30][25] , \read_value_mux[30][24] ,
         \read_value_mux[30][23] , \read_value_mux[30][22] ,
         \read_value_mux[30][21] , \read_value_mux[30][20] ,
         \read_value_mux[30][19] , \read_value_mux[30][18] ,
         \read_value_mux[30][17] , \read_value_mux[30][16] ,
         \read_value_mux[30][15] , \read_value_mux[30][14] ,
         \read_value_mux[30][13] , \read_value_mux[30][12] ,
         \read_value_mux[30][11] , \read_value_mux[30][10] ,
         \read_value_mux[30][9] , \read_value_mux[30][8] ,
         \read_value_mux[30][7] , \read_value_mux[30][6] ,
         \read_value_mux[30][5] , \read_value_mux[30][4] ,
         \read_value_mux[30][3] , \read_value_mux[30][2] ,
         \read_value_mux[30][1] , \read_value_mux[30][0] ,
         \read_value_mux[29][31] , \read_value_mux[29][30] ,
         \read_value_mux[29][29] , \read_value_mux[29][28] ,
         \read_value_mux[29][27] , \read_value_mux[29][26] ,
         \read_value_mux[29][25] , \read_value_mux[29][24] ,
         \read_value_mux[29][23] , \read_value_mux[29][22] ,
         \read_value_mux[29][21] , \read_value_mux[29][20] ,
         \read_value_mux[29][19] , \read_value_mux[29][18] ,
         \read_value_mux[29][17] , \read_value_mux[29][16] ,
         \read_value_mux[29][15] , \read_value_mux[29][14] ,
         \read_value_mux[29][13] , \read_value_mux[29][12] ,
         \read_value_mux[29][11] , \read_value_mux[29][10] ,
         \read_value_mux[29][9] , \read_value_mux[29][8] ,
         \read_value_mux[29][7] , \read_value_mux[29][6] ,
         \read_value_mux[29][5] , \read_value_mux[29][4] ,
         \read_value_mux[29][3] , \read_value_mux[29][2] ,
         \read_value_mux[29][1] , \read_value_mux[29][0] ,
         \read_value_mux[28][31] , \read_value_mux[28][30] ,
         \read_value_mux[28][29] , \read_value_mux[28][28] ,
         \read_value_mux[28][27] , \read_value_mux[28][26] ,
         \read_value_mux[28][25] , \read_value_mux[28][24] ,
         \read_value_mux[28][23] , \read_value_mux[28][22] ,
         \read_value_mux[28][21] , \read_value_mux[28][20] ,
         \read_value_mux[28][19] , \read_value_mux[28][18] ,
         \read_value_mux[28][17] , \read_value_mux[28][16] ,
         \read_value_mux[28][15] , \read_value_mux[28][14] ,
         \read_value_mux[28][13] , \read_value_mux[28][12] ,
         \read_value_mux[28][11] , \read_value_mux[28][10] ,
         \read_value_mux[28][9] , \read_value_mux[28][8] ,
         \read_value_mux[28][7] , \read_value_mux[28][6] ,
         \read_value_mux[28][5] , \read_value_mux[28][4] ,
         \read_value_mux[28][3] , \read_value_mux[28][2] ,
         \read_value_mux[28][1] , \read_value_mux[28][0] ,
         \read_value_mux[27][31] , \read_value_mux[27][30] ,
         \read_value_mux[27][29] , \read_value_mux[27][28] ,
         \read_value_mux[27][27] , \read_value_mux[27][26] ,
         \read_value_mux[27][25] , \read_value_mux[27][24] ,
         \read_value_mux[27][23] , \read_value_mux[27][22] ,
         \read_value_mux[27][21] , \read_value_mux[27][20] ,
         \read_value_mux[27][19] , \read_value_mux[27][18] ,
         \read_value_mux[27][17] , \read_value_mux[27][16] ,
         \read_value_mux[27][15] , \read_value_mux[27][14] ,
         \read_value_mux[27][13] , \read_value_mux[27][12] ,
         \read_value_mux[27][11] , \read_value_mux[27][10] ,
         \read_value_mux[27][9] , \read_value_mux[27][8] ,
         \read_value_mux[27][7] , \read_value_mux[27][6] ,
         \read_value_mux[27][5] , \read_value_mux[27][4] ,
         \read_value_mux[27][3] , \read_value_mux[27][2] ,
         \read_value_mux[27][1] , \read_value_mux[27][0] ,
         \read_value_mux[26][31] , \read_value_mux[26][30] ,
         \read_value_mux[26][29] , \read_value_mux[26][28] ,
         \read_value_mux[26][27] , \read_value_mux[26][26] ,
         \read_value_mux[26][25] , \read_value_mux[26][24] ,
         \read_value_mux[26][23] , \read_value_mux[26][22] ,
         \read_value_mux[26][21] , \read_value_mux[26][20] ,
         \read_value_mux[26][19] , \read_value_mux[26][18] ,
         \read_value_mux[26][17] , \read_value_mux[26][16] ,
         \read_value_mux[26][15] , \read_value_mux[26][14] ,
         \read_value_mux[26][13] , \read_value_mux[26][12] ,
         \read_value_mux[26][11] , \read_value_mux[26][10] ,
         \read_value_mux[26][9] , \read_value_mux[26][8] ,
         \read_value_mux[26][7] , \read_value_mux[26][6] ,
         \read_value_mux[26][5] , \read_value_mux[26][4] ,
         \read_value_mux[26][3] , \read_value_mux[26][2] ,
         \read_value_mux[26][1] , \read_value_mux[26][0] ,
         \read_value_mux[25][31] , \read_value_mux[25][30] ,
         \read_value_mux[25][29] , \read_value_mux[25][28] ,
         \read_value_mux[25][27] , \read_value_mux[25][26] ,
         \read_value_mux[25][25] , \read_value_mux[25][24] ,
         \read_value_mux[25][23] , \read_value_mux[25][22] ,
         \read_value_mux[25][21] , \read_value_mux[25][20] ,
         \read_value_mux[25][19] , \read_value_mux[25][18] ,
         \read_value_mux[25][17] , \read_value_mux[25][16] ,
         \read_value_mux[25][15] , \read_value_mux[25][14] ,
         \read_value_mux[25][13] , \read_value_mux[25][12] ,
         \read_value_mux[25][11] , \read_value_mux[25][10] ,
         \read_value_mux[25][9] , \read_value_mux[25][8] ,
         \read_value_mux[25][7] , \read_value_mux[25][6] ,
         \read_value_mux[25][5] , \read_value_mux[25][4] ,
         \read_value_mux[25][3] , \read_value_mux[25][2] ,
         \read_value_mux[25][1] , \read_value_mux[25][0] ,
         \read_value_mux[24][31] , \read_value_mux[24][30] ,
         \read_value_mux[24][29] , \read_value_mux[24][28] ,
         \read_value_mux[24][27] , \read_value_mux[24][26] ,
         \read_value_mux[24][25] , \read_value_mux[24][24] ,
         \read_value_mux[24][23] , \read_value_mux[24][22] ,
         \read_value_mux[24][21] , \read_value_mux[24][20] ,
         \read_value_mux[24][19] , \read_value_mux[24][18] ,
         \read_value_mux[24][17] , \read_value_mux[24][16] ,
         \read_value_mux[24][15] , \read_value_mux[24][14] ,
         \read_value_mux[24][13] , \read_value_mux[24][12] ,
         \read_value_mux[24][11] , \read_value_mux[24][10] ,
         \read_value_mux[24][9] , \read_value_mux[24][8] ,
         \read_value_mux[24][7] , \read_value_mux[24][6] ,
         \read_value_mux[24][5] , \read_value_mux[24][4] ,
         \read_value_mux[24][3] , \read_value_mux[24][2] ,
         \read_value_mux[24][1] , \read_value_mux[24][0] ,
         \read_value_mux[23][31] , \read_value_mux[23][30] ,
         \read_value_mux[23][29] , \read_value_mux[23][28] ,
         \read_value_mux[23][27] , \read_value_mux[23][26] ,
         \read_value_mux[23][25] , \read_value_mux[23][24] ,
         \read_value_mux[23][23] , \read_value_mux[23][22] ,
         \read_value_mux[23][21] , \read_value_mux[23][20] ,
         \read_value_mux[23][19] , \read_value_mux[23][18] ,
         \read_value_mux[23][17] , \read_value_mux[23][16] ,
         \read_value_mux[23][15] , \read_value_mux[23][14] ,
         \read_value_mux[23][13] , \read_value_mux[23][12] ,
         \read_value_mux[23][11] , \read_value_mux[23][10] ,
         \read_value_mux[23][9] , \read_value_mux[23][8] ,
         \read_value_mux[23][7] , \read_value_mux[23][6] ,
         \read_value_mux[23][5] , \read_value_mux[23][4] ,
         \read_value_mux[23][3] , \read_value_mux[23][2] ,
         \read_value_mux[23][1] , \read_value_mux[23][0] ,
         \read_value_mux[22][31] , \read_value_mux[22][30] ,
         \read_value_mux[22][29] , \read_value_mux[22][28] ,
         \read_value_mux[22][27] , \read_value_mux[22][26] ,
         \read_value_mux[22][25] , \read_value_mux[22][24] ,
         \read_value_mux[22][23] , \read_value_mux[22][22] ,
         \read_value_mux[22][21] , \read_value_mux[22][20] ,
         \read_value_mux[22][19] , \read_value_mux[22][18] ,
         \read_value_mux[22][17] , \read_value_mux[22][16] ,
         \read_value_mux[22][15] , \read_value_mux[22][14] ,
         \read_value_mux[22][13] , \read_value_mux[22][12] ,
         \read_value_mux[22][11] , \read_value_mux[22][10] ,
         \read_value_mux[22][9] , \read_value_mux[22][8] ,
         \read_value_mux[22][7] , \read_value_mux[22][6] ,
         \read_value_mux[22][5] , \read_value_mux[22][4] ,
         \read_value_mux[22][3] , \read_value_mux[22][2] ,
         \read_value_mux[22][1] , \read_value_mux[22][0] ,
         \read_value_mux[21][31] , \read_value_mux[21][30] ,
         \read_value_mux[21][29] , \read_value_mux[21][28] ,
         \read_value_mux[21][27] , \read_value_mux[21][26] ,
         \read_value_mux[21][25] , \read_value_mux[21][24] ,
         \read_value_mux[21][23] , \read_value_mux[21][22] ,
         \read_value_mux[21][21] , \read_value_mux[21][20] ,
         \read_value_mux[21][19] , \read_value_mux[21][18] ,
         \read_value_mux[21][17] , \read_value_mux[21][16] ,
         \read_value_mux[21][15] , \read_value_mux[21][14] ,
         \read_value_mux[21][13] , \read_value_mux[21][12] ,
         \read_value_mux[21][11] , \read_value_mux[21][10] ,
         \read_value_mux[21][9] , \read_value_mux[21][8] ,
         \read_value_mux[21][7] , \read_value_mux[21][6] ,
         \read_value_mux[21][5] , \read_value_mux[21][4] ,
         \read_value_mux[21][3] , \read_value_mux[21][2] ,
         \read_value_mux[21][1] , \read_value_mux[21][0] ,
         \read_value_mux[20][31] , \read_value_mux[20][30] ,
         \read_value_mux[20][29] , \read_value_mux[20][28] ,
         \read_value_mux[20][27] , \read_value_mux[20][26] ,
         \read_value_mux[20][25] , \read_value_mux[20][24] ,
         \read_value_mux[20][23] , \read_value_mux[20][22] ,
         \read_value_mux[20][21] , \read_value_mux[20][20] ,
         \read_value_mux[20][19] , \read_value_mux[20][18] ,
         \read_value_mux[20][17] , \read_value_mux[20][16] ,
         \read_value_mux[20][15] , \read_value_mux[20][14] ,
         \read_value_mux[20][13] , \read_value_mux[20][12] ,
         \read_value_mux[20][11] , \read_value_mux[20][10] ,
         \read_value_mux[20][9] , \read_value_mux[20][8] ,
         \read_value_mux[20][7] , \read_value_mux[20][6] ,
         \read_value_mux[20][5] , \read_value_mux[20][4] ,
         \read_value_mux[20][3] , \read_value_mux[20][2] ,
         \read_value_mux[20][1] , \read_value_mux[20][0] ,
         \read_value_mux[19][31] , \read_value_mux[19][30] ,
         \read_value_mux[19][29] , \read_value_mux[19][28] ,
         \read_value_mux[19][27] , \read_value_mux[19][26] ,
         \read_value_mux[19][25] , \read_value_mux[19][24] ,
         \read_value_mux[19][23] , \read_value_mux[19][22] ,
         \read_value_mux[19][21] , \read_value_mux[19][20] ,
         \read_value_mux[19][19] , \read_value_mux[19][18] ,
         \read_value_mux[19][17] , \read_value_mux[19][16] ,
         \read_value_mux[19][15] , \read_value_mux[19][14] ,
         \read_value_mux[19][13] , \read_value_mux[19][12] ,
         \read_value_mux[19][11] , \read_value_mux[19][10] ,
         \read_value_mux[19][9] , \read_value_mux[19][8] ,
         \read_value_mux[19][7] , \read_value_mux[19][6] ,
         \read_value_mux[19][5] , \read_value_mux[19][4] ,
         \read_value_mux[19][3] , \read_value_mux[19][2] ,
         \read_value_mux[19][1] , \read_value_mux[19][0] ,
         \read_value_mux[18][31] , \read_value_mux[18][30] ,
         \read_value_mux[18][29] , \read_value_mux[18][28] ,
         \read_value_mux[18][27] , \read_value_mux[18][26] ,
         \read_value_mux[18][25] , \read_value_mux[18][24] ,
         \read_value_mux[18][23] , \read_value_mux[18][22] ,
         \read_value_mux[18][21] , \read_value_mux[18][20] ,
         \read_value_mux[18][19] , \read_value_mux[18][18] ,
         \read_value_mux[18][17] , \read_value_mux[18][16] ,
         \read_value_mux[18][15] , \read_value_mux[18][14] ,
         \read_value_mux[18][13] , \read_value_mux[18][12] ,
         \read_value_mux[18][11] , \read_value_mux[18][10] ,
         \read_value_mux[18][9] , \read_value_mux[18][8] ,
         \read_value_mux[18][7] , \read_value_mux[18][6] ,
         \read_value_mux[18][5] , \read_value_mux[18][4] ,
         \read_value_mux[18][3] , \read_value_mux[18][2] ,
         \read_value_mux[18][1] , \read_value_mux[18][0] ,
         \read_value_mux[17][31] , \read_value_mux[17][30] ,
         \read_value_mux[17][29] , \read_value_mux[17][28] ,
         \read_value_mux[17][27] , \read_value_mux[17][26] ,
         \read_value_mux[17][25] , \read_value_mux[17][24] ,
         \read_value_mux[17][23] , \read_value_mux[17][22] ,
         \read_value_mux[17][21] , \read_value_mux[17][20] ,
         \read_value_mux[17][19] , \read_value_mux[17][18] ,
         \read_value_mux[17][17] , \read_value_mux[17][16] ,
         \read_value_mux[17][15] , \read_value_mux[17][14] ,
         \read_value_mux[17][13] , \read_value_mux[17][12] ,
         \read_value_mux[17][11] , \read_value_mux[17][10] ,
         \read_value_mux[17][9] , \read_value_mux[17][8] ,
         \read_value_mux[17][7] , \read_value_mux[17][6] ,
         \read_value_mux[17][5] , \read_value_mux[17][4] ,
         \read_value_mux[17][3] , \read_value_mux[17][2] ,
         \read_value_mux[17][1] , \read_value_mux[17][0] ,
         \read_value_mux[16][31] , \read_value_mux[16][30] ,
         \read_value_mux[16][29] , \read_value_mux[16][28] ,
         \read_value_mux[16][27] , \read_value_mux[16][26] ,
         \read_value_mux[16][25] , \read_value_mux[16][24] ,
         \read_value_mux[16][23] , \read_value_mux[16][22] ,
         \read_value_mux[16][21] , \read_value_mux[16][20] ,
         \read_value_mux[16][19] , \read_value_mux[16][18] ,
         \read_value_mux[16][17] , \read_value_mux[16][16] ,
         \read_value_mux[16][15] , \read_value_mux[16][14] ,
         \read_value_mux[16][13] , \read_value_mux[16][12] ,
         \read_value_mux[16][11] , \read_value_mux[16][10] ,
         \read_value_mux[16][9] , \read_value_mux[16][8] ,
         \read_value_mux[16][7] , \read_value_mux[16][6] ,
         \read_value_mux[16][5] , \read_value_mux[16][4] ,
         \read_value_mux[16][3] , \read_value_mux[16][2] ,
         \read_value_mux[16][1] , \read_value_mux[16][0] ,
         \read_value_mux[15][31] , \read_value_mux[15][30] ,
         \read_value_mux[15][29] , \read_value_mux[15][28] ,
         \read_value_mux[15][27] , \read_value_mux[15][26] ,
         \read_value_mux[15][25] , \read_value_mux[15][24] ,
         \read_value_mux[15][23] , \read_value_mux[15][22] ,
         \read_value_mux[15][21] , \read_value_mux[15][20] ,
         \read_value_mux[15][19] , \read_value_mux[15][18] ,
         \read_value_mux[15][17] , \read_value_mux[15][16] ,
         \read_value_mux[15][15] , \read_value_mux[15][14] ,
         \read_value_mux[15][13] , \read_value_mux[15][12] ,
         \read_value_mux[15][11] , \read_value_mux[15][10] ,
         \read_value_mux[15][9] , \read_value_mux[15][8] ,
         \read_value_mux[15][7] , \read_value_mux[15][6] ,
         \read_value_mux[15][5] , \read_value_mux[15][4] ,
         \read_value_mux[15][3] , \read_value_mux[15][2] ,
         \read_value_mux[15][1] , \read_value_mux[15][0] ,
         \read_value_mux[14][31] , \read_value_mux[14][30] ,
         \read_value_mux[14][29] , \read_value_mux[14][28] ,
         \read_value_mux[14][27] , \read_value_mux[14][26] ,
         \read_value_mux[14][25] , \read_value_mux[14][24] ,
         \read_value_mux[14][23] , \read_value_mux[14][22] ,
         \read_value_mux[14][21] , \read_value_mux[14][20] ,
         \read_value_mux[14][19] , \read_value_mux[14][18] ,
         \read_value_mux[14][17] , \read_value_mux[14][16] ,
         \read_value_mux[14][15] , \read_value_mux[14][14] ,
         \read_value_mux[14][13] , \read_value_mux[14][12] ,
         \read_value_mux[14][11] , \read_value_mux[14][10] ,
         \read_value_mux[14][9] , \read_value_mux[14][8] ,
         \read_value_mux[14][7] , \read_value_mux[14][6] ,
         \read_value_mux[14][5] , \read_value_mux[14][4] ,
         \read_value_mux[14][3] , \read_value_mux[14][2] ,
         \read_value_mux[14][1] , \read_value_mux[14][0] ,
         \read_value_mux[13][31] , \read_value_mux[13][30] ,
         \read_value_mux[13][29] , \read_value_mux[13][28] ,
         \read_value_mux[13][27] , \read_value_mux[13][26] ,
         \read_value_mux[13][25] , \read_value_mux[13][24] ,
         \read_value_mux[13][23] , \read_value_mux[13][22] ,
         \read_value_mux[13][21] , \read_value_mux[13][20] ,
         \read_value_mux[13][19] , \read_value_mux[13][18] ,
         \read_value_mux[13][17] , \read_value_mux[13][16] ,
         \read_value_mux[13][15] , \read_value_mux[13][14] ,
         \read_value_mux[13][13] , \read_value_mux[13][12] ,
         \read_value_mux[13][11] , \read_value_mux[13][10] ,
         \read_value_mux[13][9] , \read_value_mux[13][8] ,
         \read_value_mux[13][7] , \read_value_mux[13][6] ,
         \read_value_mux[13][5] , \read_value_mux[13][4] ,
         \read_value_mux[13][3] , \read_value_mux[13][2] ,
         \read_value_mux[13][1] , \read_value_mux[13][0] ,
         \read_value_mux[12][31] , \read_value_mux[12][30] ,
         \read_value_mux[12][29] , \read_value_mux[12][28] ,
         \read_value_mux[12][27] , \read_value_mux[12][26] ,
         \read_value_mux[12][25] , \read_value_mux[12][24] ,
         \read_value_mux[12][23] , \read_value_mux[12][22] ,
         \read_value_mux[12][21] , \read_value_mux[12][20] ,
         \read_value_mux[12][19] , \read_value_mux[12][18] ,
         \read_value_mux[12][17] , \read_value_mux[12][16] ,
         \read_value_mux[12][15] , \read_value_mux[12][14] ,
         \read_value_mux[12][13] , \read_value_mux[12][12] ,
         \read_value_mux[12][11] , \read_value_mux[12][10] ,
         \read_value_mux[12][9] , \read_value_mux[12][8] ,
         \read_value_mux[12][7] , \read_value_mux[12][6] ,
         \read_value_mux[12][5] , \read_value_mux[12][4] ,
         \read_value_mux[12][3] , \read_value_mux[12][2] ,
         \read_value_mux[12][1] , \read_value_mux[12][0] ,
         \read_value_mux[11][31] , \read_value_mux[11][30] ,
         \read_value_mux[11][29] , \read_value_mux[11][28] ,
         \read_value_mux[11][27] , \read_value_mux[11][26] ,
         \read_value_mux[11][25] , \read_value_mux[11][24] ,
         \read_value_mux[11][23] , \read_value_mux[11][22] ,
         \read_value_mux[11][21] , \read_value_mux[11][20] ,
         \read_value_mux[11][19] , \read_value_mux[11][18] ,
         \read_value_mux[11][17] , \read_value_mux[11][16] ,
         \read_value_mux[11][15] , \read_value_mux[11][14] ,
         \read_value_mux[11][13] , \read_value_mux[11][12] ,
         \read_value_mux[11][11] , \read_value_mux[11][10] ,
         \read_value_mux[11][9] , \read_value_mux[11][8] ,
         \read_value_mux[11][7] , \read_value_mux[11][6] ,
         \read_value_mux[11][5] , \read_value_mux[11][4] ,
         \read_value_mux[11][3] , \read_value_mux[11][2] ,
         \read_value_mux[11][1] , \read_value_mux[11][0] ,
         \read_value_mux[10][31] , \read_value_mux[10][30] ,
         \read_value_mux[10][29] , \read_value_mux[10][28] ,
         \read_value_mux[10][27] , \read_value_mux[10][26] ,
         \read_value_mux[10][25] , \read_value_mux[10][24] ,
         \read_value_mux[10][23] , \read_value_mux[10][22] ,
         \read_value_mux[10][21] , \read_value_mux[10][20] ,
         \read_value_mux[10][19] , \read_value_mux[10][18] ,
         \read_value_mux[10][17] , \read_value_mux[10][16] ,
         \read_value_mux[10][15] , \read_value_mux[10][14] ,
         \read_value_mux[10][13] , \read_value_mux[10][12] ,
         \read_value_mux[10][11] , \read_value_mux[10][10] ,
         \read_value_mux[10][9] , \read_value_mux[10][8] ,
         \read_value_mux[10][7] , \read_value_mux[10][6] ,
         \read_value_mux[10][5] , \read_value_mux[10][4] ,
         \read_value_mux[10][3] , \read_value_mux[10][2] ,
         \read_value_mux[10][1] , \read_value_mux[10][0] ,
         \read_value_mux[9][31] , \read_value_mux[9][30] ,
         \read_value_mux[9][29] , \read_value_mux[9][28] ,
         \read_value_mux[9][27] , \read_value_mux[9][26] ,
         \read_value_mux[9][25] , \read_value_mux[9][24] ,
         \read_value_mux[9][23] , \read_value_mux[9][22] ,
         \read_value_mux[9][21] , \read_value_mux[9][20] ,
         \read_value_mux[9][19] , \read_value_mux[9][18] ,
         \read_value_mux[9][17] , \read_value_mux[9][16] ,
         \read_value_mux[9][15] , \read_value_mux[9][14] ,
         \read_value_mux[9][13] , \read_value_mux[9][12] ,
         \read_value_mux[9][11] , \read_value_mux[9][10] ,
         \read_value_mux[9][9] , \read_value_mux[9][8] ,
         \read_value_mux[9][7] , \read_value_mux[9][6] ,
         \read_value_mux[9][5] , \read_value_mux[9][4] ,
         \read_value_mux[9][3] , \read_value_mux[9][2] ,
         \read_value_mux[9][1] , \read_value_mux[9][0] ,
         \read_value_mux[8][31] , \read_value_mux[8][30] ,
         \read_value_mux[8][29] , \read_value_mux[8][28] ,
         \read_value_mux[8][27] , \read_value_mux[8][26] ,
         \read_value_mux[8][25] , \read_value_mux[8][24] ,
         \read_value_mux[8][23] , \read_value_mux[8][22] ,
         \read_value_mux[8][21] , \read_value_mux[8][20] ,
         \read_value_mux[8][19] , \read_value_mux[8][18] ,
         \read_value_mux[8][17] , \read_value_mux[8][16] ,
         \read_value_mux[8][15] , \read_value_mux[8][14] ,
         \read_value_mux[8][13] , \read_value_mux[8][12] ,
         \read_value_mux[8][11] , \read_value_mux[8][10] ,
         \read_value_mux[8][9] , \read_value_mux[8][8] ,
         \read_value_mux[8][7] , \read_value_mux[8][6] ,
         \read_value_mux[8][5] , \read_value_mux[8][4] ,
         \read_value_mux[8][3] , \read_value_mux[8][2] ,
         \read_value_mux[8][1] , \read_value_mux[8][0] ,
         \read_value_mux[7][31] , \read_value_mux[7][30] ,
         \read_value_mux[7][29] , \read_value_mux[7][28] ,
         \read_value_mux[7][27] , \read_value_mux[7][26] ,
         \read_value_mux[7][25] , \read_value_mux[7][24] ,
         \read_value_mux[7][23] , \read_value_mux[7][22] ,
         \read_value_mux[7][21] , \read_value_mux[7][20] ,
         \read_value_mux[7][19] , \read_value_mux[7][18] ,
         \read_value_mux[7][17] , \read_value_mux[7][16] ,
         \read_value_mux[7][15] , \read_value_mux[7][14] ,
         \read_value_mux[7][13] , \read_value_mux[7][12] ,
         \read_value_mux[7][11] , \read_value_mux[7][10] ,
         \read_value_mux[7][9] , \read_value_mux[7][8] ,
         \read_value_mux[7][7] , \read_value_mux[7][6] ,
         \read_value_mux[7][5] , \read_value_mux[7][4] ,
         \read_value_mux[7][3] , \read_value_mux[7][2] ,
         \read_value_mux[7][1] , \read_value_mux[7][0] ,
         \read_value_mux[6][31] , \read_value_mux[6][30] ,
         \read_value_mux[6][29] , \read_value_mux[6][28] ,
         \read_value_mux[6][27] , \read_value_mux[6][26] ,
         \read_value_mux[6][25] , \read_value_mux[6][24] ,
         \read_value_mux[6][23] , \read_value_mux[6][22] ,
         \read_value_mux[6][21] , \read_value_mux[6][20] ,
         \read_value_mux[6][19] , \read_value_mux[6][18] ,
         \read_value_mux[6][17] , \read_value_mux[6][16] ,
         \read_value_mux[6][15] , \read_value_mux[6][14] ,
         \read_value_mux[6][13] , \read_value_mux[6][12] ,
         \read_value_mux[6][11] , \read_value_mux[6][10] ,
         \read_value_mux[6][9] , \read_value_mux[6][8] ,
         \read_value_mux[6][7] , \read_value_mux[6][6] ,
         \read_value_mux[6][5] , \read_value_mux[6][4] ,
         \read_value_mux[6][3] , \read_value_mux[6][2] ,
         \read_value_mux[6][1] , \read_value_mux[6][0] ,
         \read_value_mux[5][31] , \read_value_mux[5][30] ,
         \read_value_mux[5][29] , \read_value_mux[5][28] ,
         \read_value_mux[5][27] , \read_value_mux[5][26] ,
         \read_value_mux[5][25] , \read_value_mux[5][24] ,
         \read_value_mux[5][23] , \read_value_mux[5][22] ,
         \read_value_mux[5][21] , \read_value_mux[5][20] ,
         \read_value_mux[5][19] , \read_value_mux[5][18] ,
         \read_value_mux[5][17] , \read_value_mux[5][16] ,
         \read_value_mux[5][15] , \read_value_mux[5][14] ,
         \read_value_mux[5][13] , \read_value_mux[5][12] ,
         \read_value_mux[5][11] , \read_value_mux[5][10] ,
         \read_value_mux[5][9] , \read_value_mux[5][8] ,
         \read_value_mux[5][7] , \read_value_mux[5][6] ,
         \read_value_mux[5][5] , \read_value_mux[5][4] ,
         \read_value_mux[5][3] , \read_value_mux[5][2] ,
         \read_value_mux[5][1] , \read_value_mux[5][0] ,
         \read_value_mux[4][31] , \read_value_mux[4][30] ,
         \read_value_mux[4][29] , \read_value_mux[4][28] ,
         \read_value_mux[4][27] , \read_value_mux[4][26] ,
         \read_value_mux[4][25] , \read_value_mux[4][24] ,
         \read_value_mux[4][23] , \read_value_mux[4][22] ,
         \read_value_mux[4][21] , \read_value_mux[4][20] ,
         \read_value_mux[4][19] , \read_value_mux[4][18] ,
         \read_value_mux[4][17] , \read_value_mux[4][16] ,
         \read_value_mux[4][15] , \read_value_mux[4][14] ,
         \read_value_mux[4][13] , \read_value_mux[4][12] ,
         \read_value_mux[4][11] , \read_value_mux[4][10] ,
         \read_value_mux[4][9] , \read_value_mux[4][8] ,
         \read_value_mux[4][7] , \read_value_mux[4][6] ,
         \read_value_mux[4][5] , \read_value_mux[4][4] ,
         \read_value_mux[4][3] , \read_value_mux[4][2] ,
         \read_value_mux[4][1] , \read_value_mux[4][0] ,
         \read_value_mux[3][31] , \read_value_mux[3][30] ,
         \read_value_mux[3][29] , \read_value_mux[3][28] ,
         \read_value_mux[3][27] , \read_value_mux[3][26] ,
         \read_value_mux[3][25] , \read_value_mux[3][24] ,
         \read_value_mux[3][23] , \read_value_mux[3][22] ,
         \read_value_mux[3][21] , \read_value_mux[3][20] ,
         \read_value_mux[3][19] , \read_value_mux[3][18] ,
         \read_value_mux[3][17] , \read_value_mux[3][16] ,
         \read_value_mux[3][15] , \read_value_mux[3][14] ,
         \read_value_mux[3][13] , \read_value_mux[3][12] ,
         \read_value_mux[3][11] , \read_value_mux[3][10] ,
         \read_value_mux[3][9] , \read_value_mux[3][8] ,
         \read_value_mux[3][7] , \read_value_mux[3][6] ,
         \read_value_mux[3][5] , \read_value_mux[3][4] ,
         \read_value_mux[3][3] , \read_value_mux[3][2] ,
         \read_value_mux[3][1] , \read_value_mux[3][0] ,
         \read_value_mux[2][31] , \read_value_mux[2][30] ,
         \read_value_mux[2][29] , \read_value_mux[2][28] ,
         \read_value_mux[2][27] , \read_value_mux[2][26] ,
         \read_value_mux[2][25] , \read_value_mux[2][24] ,
         \read_value_mux[2][23] , \read_value_mux[2][22] ,
         \read_value_mux[2][21] , \read_value_mux[2][20] ,
         \read_value_mux[2][19] , \read_value_mux[2][18] ,
         \read_value_mux[2][17] , \read_value_mux[2][16] ,
         \read_value_mux[2][15] , \read_value_mux[2][14] ,
         \read_value_mux[2][13] , \read_value_mux[2][12] ,
         \read_value_mux[2][11] , \read_value_mux[2][10] ,
         \read_value_mux[2][9] , \read_value_mux[2][8] ,
         \read_value_mux[2][7] , \read_value_mux[2][6] ,
         \read_value_mux[2][5] , \read_value_mux[2][4] ,
         \read_value_mux[2][3] , \read_value_mux[2][2] ,
         \read_value_mux[2][1] , \read_value_mux[2][0] ,
         \read_value_mux[1][31] , \read_value_mux[1][30] ,
         \read_value_mux[1][29] , \read_value_mux[1][28] ,
         \read_value_mux[1][27] , \read_value_mux[1][26] ,
         \read_value_mux[1][25] , \read_value_mux[1][24] ,
         \read_value_mux[1][23] , \read_value_mux[1][22] ,
         \read_value_mux[1][21] , \read_value_mux[1][20] ,
         \read_value_mux[1][19] , \read_value_mux[1][18] ,
         \read_value_mux[1][17] , \read_value_mux[1][16] ,
         \read_value_mux[1][15] , \read_value_mux[1][14] ,
         \read_value_mux[1][13] , \read_value_mux[1][12] ,
         \read_value_mux[1][11] , \read_value_mux[1][10] ,
         \read_value_mux[1][9] , \read_value_mux[1][8] ,
         \read_value_mux[1][7] , \read_value_mux[1][6] ,
         \read_value_mux[1][5] , \read_value_mux[1][4] ,
         \read_value_mux[1][3] , \read_value_mux[1][2] ,
         \read_value_mux[1][1] , \read_value_mux[1][0] ,
         \read_value_mux[0][31] , \read_value_mux[0][30] ,
         \read_value_mux[0][29] , \read_value_mux[0][28] ,
         \read_value_mux[0][27] , \read_value_mux[0][26] ,
         \read_value_mux[0][25] , \read_value_mux[0][24] ,
         \read_value_mux[0][23] , \read_value_mux[0][22] ,
         \read_value_mux[0][21] , \read_value_mux[0][20] ,
         \read_value_mux[0][19] , \read_value_mux[0][18] ,
         \read_value_mux[0][17] , \read_value_mux[0][16] ,
         \read_value_mux[0][15] , \read_value_mux[0][14] ,
         \read_value_mux[0][13] , \read_value_mux[0][12] ,
         \read_value_mux[0][11] , \read_value_mux[0][10] ,
         \read_value_mux[0][9] , \read_value_mux[0][8] ,
         \read_value_mux[0][7] , \read_value_mux[0][6] ,
         \read_value_mux[0][5] , \read_value_mux[0][4] ,
         \read_value_mux[0][3] , \read_value_mux[0][2] ,
         \read_value_mux[0][1] , \read_value_mux[0][0] , n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40;
  wire   [31:0] dec_read_index;
  wire   [31:0] dec_write_index;
  wire   [31:0] search_results;
  wire   [31:0] read_results;

  cam_word_0 \words[0]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[0]), .write(write), .dec_write_index(
        dec_write_index[0]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[0]), 
        .read_results(read_results[0]), .read_value({\read_value_mux[0][31] , 
        \read_value_mux[0][30] , \read_value_mux[0][29] , 
        \read_value_mux[0][28] , \read_value_mux[0][27] , 
        \read_value_mux[0][26] , \read_value_mux[0][25] , 
        \read_value_mux[0][24] , \read_value_mux[0][23] , 
        \read_value_mux[0][22] , \read_value_mux[0][21] , 
        \read_value_mux[0][20] , \read_value_mux[0][19] , 
        \read_value_mux[0][18] , \read_value_mux[0][17] , 
        \read_value_mux[0][16] , \read_value_mux[0][15] , 
        \read_value_mux[0][14] , \read_value_mux[0][13] , 
        \read_value_mux[0][12] , \read_value_mux[0][11] , 
        \read_value_mux[0][10] , \read_value_mux[0][9] , 
        \read_value_mux[0][8] , \read_value_mux[0][7] , \read_value_mux[0][6] , 
        \read_value_mux[0][5] , \read_value_mux[0][4] , \read_value_mux[0][3] , 
        \read_value_mux[0][2] , \read_value_mux[0][1] , \read_value_mux[0][0] }) );
  cam_word_1 \words[1]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[1]), .write(write), .dec_write_index(
        dec_write_index[1]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[1]), 
        .read_results(read_results[1]), .read_value({\read_value_mux[1][31] , 
        \read_value_mux[1][30] , \read_value_mux[1][29] , 
        \read_value_mux[1][28] , \read_value_mux[1][27] , 
        \read_value_mux[1][26] , \read_value_mux[1][25] , 
        \read_value_mux[1][24] , \read_value_mux[1][23] , 
        \read_value_mux[1][22] , \read_value_mux[1][21] , 
        \read_value_mux[1][20] , \read_value_mux[1][19] , 
        \read_value_mux[1][18] , \read_value_mux[1][17] , 
        \read_value_mux[1][16] , \read_value_mux[1][15] , 
        \read_value_mux[1][14] , \read_value_mux[1][13] , 
        \read_value_mux[1][12] , \read_value_mux[1][11] , 
        \read_value_mux[1][10] , \read_value_mux[1][9] , 
        \read_value_mux[1][8] , \read_value_mux[1][7] , \read_value_mux[1][6] , 
        \read_value_mux[1][5] , \read_value_mux[1][4] , \read_value_mux[1][3] , 
        \read_value_mux[1][2] , \read_value_mux[1][1] , \read_value_mux[1][0] }) );
  cam_word_2 \words[2]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[2]), .write(write), .dec_write_index(
        dec_write_index[2]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[2]), 
        .read_results(read_results[2]), .read_value({\read_value_mux[2][31] , 
        \read_value_mux[2][30] , \read_value_mux[2][29] , 
        \read_value_mux[2][28] , \read_value_mux[2][27] , 
        \read_value_mux[2][26] , \read_value_mux[2][25] , 
        \read_value_mux[2][24] , \read_value_mux[2][23] , 
        \read_value_mux[2][22] , \read_value_mux[2][21] , 
        \read_value_mux[2][20] , \read_value_mux[2][19] , 
        \read_value_mux[2][18] , \read_value_mux[2][17] , 
        \read_value_mux[2][16] , \read_value_mux[2][15] , 
        \read_value_mux[2][14] , \read_value_mux[2][13] , 
        \read_value_mux[2][12] , \read_value_mux[2][11] , 
        \read_value_mux[2][10] , \read_value_mux[2][9] , 
        \read_value_mux[2][8] , \read_value_mux[2][7] , \read_value_mux[2][6] , 
        \read_value_mux[2][5] , \read_value_mux[2][4] , \read_value_mux[2][3] , 
        \read_value_mux[2][2] , \read_value_mux[2][1] , \read_value_mux[2][0] }) );
  cam_word_3 \words[3]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[3]), .write(write), .dec_write_index(
        dec_write_index[3]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[3]), 
        .read_results(read_results[3]), .read_value({\read_value_mux[3][31] , 
        \read_value_mux[3][30] , \read_value_mux[3][29] , 
        \read_value_mux[3][28] , \read_value_mux[3][27] , 
        \read_value_mux[3][26] , \read_value_mux[3][25] , 
        \read_value_mux[3][24] , \read_value_mux[3][23] , 
        \read_value_mux[3][22] , \read_value_mux[3][21] , 
        \read_value_mux[3][20] , \read_value_mux[3][19] , 
        \read_value_mux[3][18] , \read_value_mux[3][17] , 
        \read_value_mux[3][16] , \read_value_mux[3][15] , 
        \read_value_mux[3][14] , \read_value_mux[3][13] , 
        \read_value_mux[3][12] , \read_value_mux[3][11] , 
        \read_value_mux[3][10] , \read_value_mux[3][9] , 
        \read_value_mux[3][8] , \read_value_mux[3][7] , \read_value_mux[3][6] , 
        \read_value_mux[3][5] , \read_value_mux[3][4] , \read_value_mux[3][3] , 
        \read_value_mux[3][2] , \read_value_mux[3][1] , \read_value_mux[3][0] }) );
  cam_word_4 \words[4]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[4]), .write(write), .dec_write_index(
        dec_write_index[4]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[4]), 
        .read_results(read_results[4]), .read_value({\read_value_mux[4][31] , 
        \read_value_mux[4][30] , \read_value_mux[4][29] , 
        \read_value_mux[4][28] , \read_value_mux[4][27] , 
        \read_value_mux[4][26] , \read_value_mux[4][25] , 
        \read_value_mux[4][24] , \read_value_mux[4][23] , 
        \read_value_mux[4][22] , \read_value_mux[4][21] , 
        \read_value_mux[4][20] , \read_value_mux[4][19] , 
        \read_value_mux[4][18] , \read_value_mux[4][17] , 
        \read_value_mux[4][16] , \read_value_mux[4][15] , 
        \read_value_mux[4][14] , \read_value_mux[4][13] , 
        \read_value_mux[4][12] , \read_value_mux[4][11] , 
        \read_value_mux[4][10] , \read_value_mux[4][9] , 
        \read_value_mux[4][8] , \read_value_mux[4][7] , \read_value_mux[4][6] , 
        \read_value_mux[4][5] , \read_value_mux[4][4] , \read_value_mux[4][3] , 
        \read_value_mux[4][2] , \read_value_mux[4][1] , \read_value_mux[4][0] }) );
  cam_word_5 \words[5]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[5]), .write(write), .dec_write_index(
        dec_write_index[5]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[5]), 
        .read_results(read_results[5]), .read_value({\read_value_mux[5][31] , 
        \read_value_mux[5][30] , \read_value_mux[5][29] , 
        \read_value_mux[5][28] , \read_value_mux[5][27] , 
        \read_value_mux[5][26] , \read_value_mux[5][25] , 
        \read_value_mux[5][24] , \read_value_mux[5][23] , 
        \read_value_mux[5][22] , \read_value_mux[5][21] , 
        \read_value_mux[5][20] , \read_value_mux[5][19] , 
        \read_value_mux[5][18] , \read_value_mux[5][17] , 
        \read_value_mux[5][16] , \read_value_mux[5][15] , 
        \read_value_mux[5][14] , \read_value_mux[5][13] , 
        \read_value_mux[5][12] , \read_value_mux[5][11] , 
        \read_value_mux[5][10] , \read_value_mux[5][9] , 
        \read_value_mux[5][8] , \read_value_mux[5][7] , \read_value_mux[5][6] , 
        \read_value_mux[5][5] , \read_value_mux[5][4] , \read_value_mux[5][3] , 
        \read_value_mux[5][2] , \read_value_mux[5][1] , \read_value_mux[5][0] }) );
  cam_word_6 \words[6]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[6]), .write(write), .dec_write_index(
        dec_write_index[6]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[6]), 
        .read_results(read_results[6]), .read_value({\read_value_mux[6][31] , 
        \read_value_mux[6][30] , \read_value_mux[6][29] , 
        \read_value_mux[6][28] , \read_value_mux[6][27] , 
        \read_value_mux[6][26] , \read_value_mux[6][25] , 
        \read_value_mux[6][24] , \read_value_mux[6][23] , 
        \read_value_mux[6][22] , \read_value_mux[6][21] , 
        \read_value_mux[6][20] , \read_value_mux[6][19] , 
        \read_value_mux[6][18] , \read_value_mux[6][17] , 
        \read_value_mux[6][16] , \read_value_mux[6][15] , 
        \read_value_mux[6][14] , \read_value_mux[6][13] , 
        \read_value_mux[6][12] , \read_value_mux[6][11] , 
        \read_value_mux[6][10] , \read_value_mux[6][9] , 
        \read_value_mux[6][8] , \read_value_mux[6][7] , \read_value_mux[6][6] , 
        \read_value_mux[6][5] , \read_value_mux[6][4] , \read_value_mux[6][3] , 
        \read_value_mux[6][2] , \read_value_mux[6][1] , \read_value_mux[6][0] }) );
  cam_word_7 \words[7]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[7]), .write(write), .dec_write_index(
        dec_write_index[7]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[7]), 
        .read_results(read_results[7]), .read_value({\read_value_mux[7][31] , 
        \read_value_mux[7][30] , \read_value_mux[7][29] , 
        \read_value_mux[7][28] , \read_value_mux[7][27] , 
        \read_value_mux[7][26] , \read_value_mux[7][25] , 
        \read_value_mux[7][24] , \read_value_mux[7][23] , 
        \read_value_mux[7][22] , \read_value_mux[7][21] , 
        \read_value_mux[7][20] , \read_value_mux[7][19] , 
        \read_value_mux[7][18] , \read_value_mux[7][17] , 
        \read_value_mux[7][16] , \read_value_mux[7][15] , 
        \read_value_mux[7][14] , \read_value_mux[7][13] , 
        \read_value_mux[7][12] , \read_value_mux[7][11] , 
        \read_value_mux[7][10] , \read_value_mux[7][9] , 
        \read_value_mux[7][8] , \read_value_mux[7][7] , \read_value_mux[7][6] , 
        \read_value_mux[7][5] , \read_value_mux[7][4] , \read_value_mux[7][3] , 
        \read_value_mux[7][2] , \read_value_mux[7][1] , \read_value_mux[7][0] }) );
  cam_word_8 \words[8]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[8]), .write(write), .dec_write_index(
        dec_write_index[8]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[8]), 
        .read_results(read_results[8]), .read_value({\read_value_mux[8][31] , 
        \read_value_mux[8][30] , \read_value_mux[8][29] , 
        \read_value_mux[8][28] , \read_value_mux[8][27] , 
        \read_value_mux[8][26] , \read_value_mux[8][25] , 
        \read_value_mux[8][24] , \read_value_mux[8][23] , 
        \read_value_mux[8][22] , \read_value_mux[8][21] , 
        \read_value_mux[8][20] , \read_value_mux[8][19] , 
        \read_value_mux[8][18] , \read_value_mux[8][17] , 
        \read_value_mux[8][16] , \read_value_mux[8][15] , 
        \read_value_mux[8][14] , \read_value_mux[8][13] , 
        \read_value_mux[8][12] , \read_value_mux[8][11] , 
        \read_value_mux[8][10] , \read_value_mux[8][9] , 
        \read_value_mux[8][8] , \read_value_mux[8][7] , \read_value_mux[8][6] , 
        \read_value_mux[8][5] , \read_value_mux[8][4] , \read_value_mux[8][3] , 
        \read_value_mux[8][2] , \read_value_mux[8][1] , \read_value_mux[8][0] }) );
  cam_word_9 \words[9]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[9]), .write(write), .dec_write_index(
        dec_write_index[9]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[9]), 
        .read_results(read_results[9]), .read_value({\read_value_mux[9][31] , 
        \read_value_mux[9][30] , \read_value_mux[9][29] , 
        \read_value_mux[9][28] , \read_value_mux[9][27] , 
        \read_value_mux[9][26] , \read_value_mux[9][25] , 
        \read_value_mux[9][24] , \read_value_mux[9][23] , 
        \read_value_mux[9][22] , \read_value_mux[9][21] , 
        \read_value_mux[9][20] , \read_value_mux[9][19] , 
        \read_value_mux[9][18] , \read_value_mux[9][17] , 
        \read_value_mux[9][16] , \read_value_mux[9][15] , 
        \read_value_mux[9][14] , \read_value_mux[9][13] , 
        \read_value_mux[9][12] , \read_value_mux[9][11] , 
        \read_value_mux[9][10] , \read_value_mux[9][9] , 
        \read_value_mux[9][8] , \read_value_mux[9][7] , \read_value_mux[9][6] , 
        \read_value_mux[9][5] , \read_value_mux[9][4] , \read_value_mux[9][3] , 
        \read_value_mux[9][2] , \read_value_mux[9][1] , \read_value_mux[9][0] }) );
  cam_word_10 \words[10]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[10]), .write(write), .dec_write_index(
        dec_write_index[10]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[10]), 
        .read_results(read_results[10]), .read_value({\read_value_mux[10][31] , 
        \read_value_mux[10][30] , \read_value_mux[10][29] , 
        \read_value_mux[10][28] , \read_value_mux[10][27] , 
        \read_value_mux[10][26] , \read_value_mux[10][25] , 
        \read_value_mux[10][24] , \read_value_mux[10][23] , 
        \read_value_mux[10][22] , \read_value_mux[10][21] , 
        \read_value_mux[10][20] , \read_value_mux[10][19] , 
        \read_value_mux[10][18] , \read_value_mux[10][17] , 
        \read_value_mux[10][16] , \read_value_mux[10][15] , 
        \read_value_mux[10][14] , \read_value_mux[10][13] , 
        \read_value_mux[10][12] , \read_value_mux[10][11] , 
        \read_value_mux[10][10] , \read_value_mux[10][9] , 
        \read_value_mux[10][8] , \read_value_mux[10][7] , 
        \read_value_mux[10][6] , \read_value_mux[10][5] , 
        \read_value_mux[10][4] , \read_value_mux[10][3] , 
        \read_value_mux[10][2] , \read_value_mux[10][1] , 
        \read_value_mux[10][0] }) );
  cam_word_11 \words[11]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[11]), .write(write), .dec_write_index(
        dec_write_index[11]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[11]), 
        .read_results(read_results[11]), .read_value({\read_value_mux[11][31] , 
        \read_value_mux[11][30] , \read_value_mux[11][29] , 
        \read_value_mux[11][28] , \read_value_mux[11][27] , 
        \read_value_mux[11][26] , \read_value_mux[11][25] , 
        \read_value_mux[11][24] , \read_value_mux[11][23] , 
        \read_value_mux[11][22] , \read_value_mux[11][21] , 
        \read_value_mux[11][20] , \read_value_mux[11][19] , 
        \read_value_mux[11][18] , \read_value_mux[11][17] , 
        \read_value_mux[11][16] , \read_value_mux[11][15] , 
        \read_value_mux[11][14] , \read_value_mux[11][13] , 
        \read_value_mux[11][12] , \read_value_mux[11][11] , 
        \read_value_mux[11][10] , \read_value_mux[11][9] , 
        \read_value_mux[11][8] , \read_value_mux[11][7] , 
        \read_value_mux[11][6] , \read_value_mux[11][5] , 
        \read_value_mux[11][4] , \read_value_mux[11][3] , 
        \read_value_mux[11][2] , \read_value_mux[11][1] , 
        \read_value_mux[11][0] }) );
  cam_word_12 \words[12]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[12]), .write(write), .dec_write_index(
        dec_write_index[12]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[12]), 
        .read_results(read_results[12]), .read_value({\read_value_mux[12][31] , 
        \read_value_mux[12][30] , \read_value_mux[12][29] , 
        \read_value_mux[12][28] , \read_value_mux[12][27] , 
        \read_value_mux[12][26] , \read_value_mux[12][25] , 
        \read_value_mux[12][24] , \read_value_mux[12][23] , 
        \read_value_mux[12][22] , \read_value_mux[12][21] , 
        \read_value_mux[12][20] , \read_value_mux[12][19] , 
        \read_value_mux[12][18] , \read_value_mux[12][17] , 
        \read_value_mux[12][16] , \read_value_mux[12][15] , 
        \read_value_mux[12][14] , \read_value_mux[12][13] , 
        \read_value_mux[12][12] , \read_value_mux[12][11] , 
        \read_value_mux[12][10] , \read_value_mux[12][9] , 
        \read_value_mux[12][8] , \read_value_mux[12][7] , 
        \read_value_mux[12][6] , \read_value_mux[12][5] , 
        \read_value_mux[12][4] , \read_value_mux[12][3] , 
        \read_value_mux[12][2] , \read_value_mux[12][1] , 
        \read_value_mux[12][0] }) );
  cam_word_13 \words[13]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[13]), .write(write), .dec_write_index(
        dec_write_index[13]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[13]), 
        .read_results(read_results[13]), .read_value({\read_value_mux[13][31] , 
        \read_value_mux[13][30] , \read_value_mux[13][29] , 
        \read_value_mux[13][28] , \read_value_mux[13][27] , 
        \read_value_mux[13][26] , \read_value_mux[13][25] , 
        \read_value_mux[13][24] , \read_value_mux[13][23] , 
        \read_value_mux[13][22] , \read_value_mux[13][21] , 
        \read_value_mux[13][20] , \read_value_mux[13][19] , 
        \read_value_mux[13][18] , \read_value_mux[13][17] , 
        \read_value_mux[13][16] , \read_value_mux[13][15] , 
        \read_value_mux[13][14] , \read_value_mux[13][13] , 
        \read_value_mux[13][12] , \read_value_mux[13][11] , 
        \read_value_mux[13][10] , \read_value_mux[13][9] , 
        \read_value_mux[13][8] , \read_value_mux[13][7] , 
        \read_value_mux[13][6] , \read_value_mux[13][5] , 
        \read_value_mux[13][4] , \read_value_mux[13][3] , 
        \read_value_mux[13][2] , \read_value_mux[13][1] , 
        \read_value_mux[13][0] }) );
  cam_word_14 \words[14]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[14]), .write(write), .dec_write_index(
        dec_write_index[14]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[14]), 
        .read_results(read_results[14]), .read_value({\read_value_mux[14][31] , 
        \read_value_mux[14][30] , \read_value_mux[14][29] , 
        \read_value_mux[14][28] , \read_value_mux[14][27] , 
        \read_value_mux[14][26] , \read_value_mux[14][25] , 
        \read_value_mux[14][24] , \read_value_mux[14][23] , 
        \read_value_mux[14][22] , \read_value_mux[14][21] , 
        \read_value_mux[14][20] , \read_value_mux[14][19] , 
        \read_value_mux[14][18] , \read_value_mux[14][17] , 
        \read_value_mux[14][16] , \read_value_mux[14][15] , 
        \read_value_mux[14][14] , \read_value_mux[14][13] , 
        \read_value_mux[14][12] , \read_value_mux[14][11] , 
        \read_value_mux[14][10] , \read_value_mux[14][9] , 
        \read_value_mux[14][8] , \read_value_mux[14][7] , 
        \read_value_mux[14][6] , \read_value_mux[14][5] , 
        \read_value_mux[14][4] , \read_value_mux[14][3] , 
        \read_value_mux[14][2] , \read_value_mux[14][1] , 
        \read_value_mux[14][0] }) );
  cam_word_15 \words[15]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[15]), .write(write), .dec_write_index(
        dec_write_index[15]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[15]), 
        .read_results(read_results[15]), .read_value({\read_value_mux[15][31] , 
        \read_value_mux[15][30] , \read_value_mux[15][29] , 
        \read_value_mux[15][28] , \read_value_mux[15][27] , 
        \read_value_mux[15][26] , \read_value_mux[15][25] , 
        \read_value_mux[15][24] , \read_value_mux[15][23] , 
        \read_value_mux[15][22] , \read_value_mux[15][21] , 
        \read_value_mux[15][20] , \read_value_mux[15][19] , 
        \read_value_mux[15][18] , \read_value_mux[15][17] , 
        \read_value_mux[15][16] , \read_value_mux[15][15] , 
        \read_value_mux[15][14] , \read_value_mux[15][13] , 
        \read_value_mux[15][12] , \read_value_mux[15][11] , 
        \read_value_mux[15][10] , \read_value_mux[15][9] , 
        \read_value_mux[15][8] , \read_value_mux[15][7] , 
        \read_value_mux[15][6] , \read_value_mux[15][5] , 
        \read_value_mux[15][4] , \read_value_mux[15][3] , 
        \read_value_mux[15][2] , \read_value_mux[15][1] , 
        \read_value_mux[15][0] }) );
  cam_word_16 \words[16]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[16]), .write(write), .dec_write_index(
        dec_write_index[16]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[16]), 
        .read_results(read_results[16]), .read_value({\read_value_mux[16][31] , 
        \read_value_mux[16][30] , \read_value_mux[16][29] , 
        \read_value_mux[16][28] , \read_value_mux[16][27] , 
        \read_value_mux[16][26] , \read_value_mux[16][25] , 
        \read_value_mux[16][24] , \read_value_mux[16][23] , 
        \read_value_mux[16][22] , \read_value_mux[16][21] , 
        \read_value_mux[16][20] , \read_value_mux[16][19] , 
        \read_value_mux[16][18] , \read_value_mux[16][17] , 
        \read_value_mux[16][16] , \read_value_mux[16][15] , 
        \read_value_mux[16][14] , \read_value_mux[16][13] , 
        \read_value_mux[16][12] , \read_value_mux[16][11] , 
        \read_value_mux[16][10] , \read_value_mux[16][9] , 
        \read_value_mux[16][8] , \read_value_mux[16][7] , 
        \read_value_mux[16][6] , \read_value_mux[16][5] , 
        \read_value_mux[16][4] , \read_value_mux[16][3] , 
        \read_value_mux[16][2] , \read_value_mux[16][1] , 
        \read_value_mux[16][0] }) );
  cam_word_17 \words[17]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[17]), .write(write), .dec_write_index(
        dec_write_index[17]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[17]), 
        .read_results(read_results[17]), .read_value({\read_value_mux[17][31] , 
        \read_value_mux[17][30] , \read_value_mux[17][29] , 
        \read_value_mux[17][28] , \read_value_mux[17][27] , 
        \read_value_mux[17][26] , \read_value_mux[17][25] , 
        \read_value_mux[17][24] , \read_value_mux[17][23] , 
        \read_value_mux[17][22] , \read_value_mux[17][21] , 
        \read_value_mux[17][20] , \read_value_mux[17][19] , 
        \read_value_mux[17][18] , \read_value_mux[17][17] , 
        \read_value_mux[17][16] , \read_value_mux[17][15] , 
        \read_value_mux[17][14] , \read_value_mux[17][13] , 
        \read_value_mux[17][12] , \read_value_mux[17][11] , 
        \read_value_mux[17][10] , \read_value_mux[17][9] , 
        \read_value_mux[17][8] , \read_value_mux[17][7] , 
        \read_value_mux[17][6] , \read_value_mux[17][5] , 
        \read_value_mux[17][4] , \read_value_mux[17][3] , 
        \read_value_mux[17][2] , \read_value_mux[17][1] , 
        \read_value_mux[17][0] }) );
  cam_word_18 \words[18]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[18]), .write(write), .dec_write_index(
        dec_write_index[18]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[18]), 
        .read_results(read_results[18]), .read_value({\read_value_mux[18][31] , 
        \read_value_mux[18][30] , \read_value_mux[18][29] , 
        \read_value_mux[18][28] , \read_value_mux[18][27] , 
        \read_value_mux[18][26] , \read_value_mux[18][25] , 
        \read_value_mux[18][24] , \read_value_mux[18][23] , 
        \read_value_mux[18][22] , \read_value_mux[18][21] , 
        \read_value_mux[18][20] , \read_value_mux[18][19] , 
        \read_value_mux[18][18] , \read_value_mux[18][17] , 
        \read_value_mux[18][16] , \read_value_mux[18][15] , 
        \read_value_mux[18][14] , \read_value_mux[18][13] , 
        \read_value_mux[18][12] , \read_value_mux[18][11] , 
        \read_value_mux[18][10] , \read_value_mux[18][9] , 
        \read_value_mux[18][8] , \read_value_mux[18][7] , 
        \read_value_mux[18][6] , \read_value_mux[18][5] , 
        \read_value_mux[18][4] , \read_value_mux[18][3] , 
        \read_value_mux[18][2] , \read_value_mux[18][1] , 
        \read_value_mux[18][0] }) );
  cam_word_19 \words[19]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[19]), .write(write), .dec_write_index(
        dec_write_index[19]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[19]), 
        .read_results(read_results[19]), .read_value({\read_value_mux[19][31] , 
        \read_value_mux[19][30] , \read_value_mux[19][29] , 
        \read_value_mux[19][28] , \read_value_mux[19][27] , 
        \read_value_mux[19][26] , \read_value_mux[19][25] , 
        \read_value_mux[19][24] , \read_value_mux[19][23] , 
        \read_value_mux[19][22] , \read_value_mux[19][21] , 
        \read_value_mux[19][20] , \read_value_mux[19][19] , 
        \read_value_mux[19][18] , \read_value_mux[19][17] , 
        \read_value_mux[19][16] , \read_value_mux[19][15] , 
        \read_value_mux[19][14] , \read_value_mux[19][13] , 
        \read_value_mux[19][12] , \read_value_mux[19][11] , 
        \read_value_mux[19][10] , \read_value_mux[19][9] , 
        \read_value_mux[19][8] , \read_value_mux[19][7] , 
        \read_value_mux[19][6] , \read_value_mux[19][5] , 
        \read_value_mux[19][4] , \read_value_mux[19][3] , 
        \read_value_mux[19][2] , \read_value_mux[19][1] , 
        \read_value_mux[19][0] }) );
  cam_word_20 \words[20]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[20]), .write(write), .dec_write_index(
        dec_write_index[20]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[20]), 
        .read_results(read_results[20]), .read_value({\read_value_mux[20][31] , 
        \read_value_mux[20][30] , \read_value_mux[20][29] , 
        \read_value_mux[20][28] , \read_value_mux[20][27] , 
        \read_value_mux[20][26] , \read_value_mux[20][25] , 
        \read_value_mux[20][24] , \read_value_mux[20][23] , 
        \read_value_mux[20][22] , \read_value_mux[20][21] , 
        \read_value_mux[20][20] , \read_value_mux[20][19] , 
        \read_value_mux[20][18] , \read_value_mux[20][17] , 
        \read_value_mux[20][16] , \read_value_mux[20][15] , 
        \read_value_mux[20][14] , \read_value_mux[20][13] , 
        \read_value_mux[20][12] , \read_value_mux[20][11] , 
        \read_value_mux[20][10] , \read_value_mux[20][9] , 
        \read_value_mux[20][8] , \read_value_mux[20][7] , 
        \read_value_mux[20][6] , \read_value_mux[20][5] , 
        \read_value_mux[20][4] , \read_value_mux[20][3] , 
        \read_value_mux[20][2] , \read_value_mux[20][1] , 
        \read_value_mux[20][0] }) );
  cam_word_21 \words[21]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[21]), .write(write), .dec_write_index(
        dec_write_index[21]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[21]), 
        .read_results(read_results[21]), .read_value({\read_value_mux[21][31] , 
        \read_value_mux[21][30] , \read_value_mux[21][29] , 
        \read_value_mux[21][28] , \read_value_mux[21][27] , 
        \read_value_mux[21][26] , \read_value_mux[21][25] , 
        \read_value_mux[21][24] , \read_value_mux[21][23] , 
        \read_value_mux[21][22] , \read_value_mux[21][21] , 
        \read_value_mux[21][20] , \read_value_mux[21][19] , 
        \read_value_mux[21][18] , \read_value_mux[21][17] , 
        \read_value_mux[21][16] , \read_value_mux[21][15] , 
        \read_value_mux[21][14] , \read_value_mux[21][13] , 
        \read_value_mux[21][12] , \read_value_mux[21][11] , 
        \read_value_mux[21][10] , \read_value_mux[21][9] , 
        \read_value_mux[21][8] , \read_value_mux[21][7] , 
        \read_value_mux[21][6] , \read_value_mux[21][5] , 
        \read_value_mux[21][4] , \read_value_mux[21][3] , 
        \read_value_mux[21][2] , \read_value_mux[21][1] , 
        \read_value_mux[21][0] }) );
  cam_word_22 \words[22]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[22]), .write(write), .dec_write_index(
        dec_write_index[22]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[22]), 
        .read_results(read_results[22]), .read_value({\read_value_mux[22][31] , 
        \read_value_mux[22][30] , \read_value_mux[22][29] , 
        \read_value_mux[22][28] , \read_value_mux[22][27] , 
        \read_value_mux[22][26] , \read_value_mux[22][25] , 
        \read_value_mux[22][24] , \read_value_mux[22][23] , 
        \read_value_mux[22][22] , \read_value_mux[22][21] , 
        \read_value_mux[22][20] , \read_value_mux[22][19] , 
        \read_value_mux[22][18] , \read_value_mux[22][17] , 
        \read_value_mux[22][16] , \read_value_mux[22][15] , 
        \read_value_mux[22][14] , \read_value_mux[22][13] , 
        \read_value_mux[22][12] , \read_value_mux[22][11] , 
        \read_value_mux[22][10] , \read_value_mux[22][9] , 
        \read_value_mux[22][8] , \read_value_mux[22][7] , 
        \read_value_mux[22][6] , \read_value_mux[22][5] , 
        \read_value_mux[22][4] , \read_value_mux[22][3] , 
        \read_value_mux[22][2] , \read_value_mux[22][1] , 
        \read_value_mux[22][0] }) );
  cam_word_23 \words[23]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[23]), .write(write), .dec_write_index(
        dec_write_index[23]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[23]), 
        .read_results(read_results[23]), .read_value({\read_value_mux[23][31] , 
        \read_value_mux[23][30] , \read_value_mux[23][29] , 
        \read_value_mux[23][28] , \read_value_mux[23][27] , 
        \read_value_mux[23][26] , \read_value_mux[23][25] , 
        \read_value_mux[23][24] , \read_value_mux[23][23] , 
        \read_value_mux[23][22] , \read_value_mux[23][21] , 
        \read_value_mux[23][20] , \read_value_mux[23][19] , 
        \read_value_mux[23][18] , \read_value_mux[23][17] , 
        \read_value_mux[23][16] , \read_value_mux[23][15] , 
        \read_value_mux[23][14] , \read_value_mux[23][13] , 
        \read_value_mux[23][12] , \read_value_mux[23][11] , 
        \read_value_mux[23][10] , \read_value_mux[23][9] , 
        \read_value_mux[23][8] , \read_value_mux[23][7] , 
        \read_value_mux[23][6] , \read_value_mux[23][5] , 
        \read_value_mux[23][4] , \read_value_mux[23][3] , 
        \read_value_mux[23][2] , \read_value_mux[23][1] , 
        \read_value_mux[23][0] }) );
  cam_word_24 \words[24]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[24]), .write(write), .dec_write_index(
        dec_write_index[24]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[24]), 
        .read_results(read_results[24]), .read_value({\read_value_mux[24][31] , 
        \read_value_mux[24][30] , \read_value_mux[24][29] , 
        \read_value_mux[24][28] , \read_value_mux[24][27] , 
        \read_value_mux[24][26] , \read_value_mux[24][25] , 
        \read_value_mux[24][24] , \read_value_mux[24][23] , 
        \read_value_mux[24][22] , \read_value_mux[24][21] , 
        \read_value_mux[24][20] , \read_value_mux[24][19] , 
        \read_value_mux[24][18] , \read_value_mux[24][17] , 
        \read_value_mux[24][16] , \read_value_mux[24][15] , 
        \read_value_mux[24][14] , \read_value_mux[24][13] , 
        \read_value_mux[24][12] , \read_value_mux[24][11] , 
        \read_value_mux[24][10] , \read_value_mux[24][9] , 
        \read_value_mux[24][8] , \read_value_mux[24][7] , 
        \read_value_mux[24][6] , \read_value_mux[24][5] , 
        \read_value_mux[24][4] , \read_value_mux[24][3] , 
        \read_value_mux[24][2] , \read_value_mux[24][1] , 
        \read_value_mux[24][0] }) );
  cam_word_25 \words[25]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[25]), .write(write), .dec_write_index(
        dec_write_index[25]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[25]), 
        .read_results(read_results[25]), .read_value({\read_value_mux[25][31] , 
        \read_value_mux[25][30] , \read_value_mux[25][29] , 
        \read_value_mux[25][28] , \read_value_mux[25][27] , 
        \read_value_mux[25][26] , \read_value_mux[25][25] , 
        \read_value_mux[25][24] , \read_value_mux[25][23] , 
        \read_value_mux[25][22] , \read_value_mux[25][21] , 
        \read_value_mux[25][20] , \read_value_mux[25][19] , 
        \read_value_mux[25][18] , \read_value_mux[25][17] , 
        \read_value_mux[25][16] , \read_value_mux[25][15] , 
        \read_value_mux[25][14] , \read_value_mux[25][13] , 
        \read_value_mux[25][12] , \read_value_mux[25][11] , 
        \read_value_mux[25][10] , \read_value_mux[25][9] , 
        \read_value_mux[25][8] , \read_value_mux[25][7] , 
        \read_value_mux[25][6] , \read_value_mux[25][5] , 
        \read_value_mux[25][4] , \read_value_mux[25][3] , 
        \read_value_mux[25][2] , \read_value_mux[25][1] , 
        \read_value_mux[25][0] }) );
  cam_word_26 \words[26]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[26]), .write(write), .dec_write_index(
        dec_write_index[26]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[26]), 
        .read_results(read_results[26]), .read_value({\read_value_mux[26][31] , 
        \read_value_mux[26][30] , \read_value_mux[26][29] , 
        \read_value_mux[26][28] , \read_value_mux[26][27] , 
        \read_value_mux[26][26] , \read_value_mux[26][25] , 
        \read_value_mux[26][24] , \read_value_mux[26][23] , 
        \read_value_mux[26][22] , \read_value_mux[26][21] , 
        \read_value_mux[26][20] , \read_value_mux[26][19] , 
        \read_value_mux[26][18] , \read_value_mux[26][17] , 
        \read_value_mux[26][16] , \read_value_mux[26][15] , 
        \read_value_mux[26][14] , \read_value_mux[26][13] , 
        \read_value_mux[26][12] , \read_value_mux[26][11] , 
        \read_value_mux[26][10] , \read_value_mux[26][9] , 
        \read_value_mux[26][8] , \read_value_mux[26][7] , 
        \read_value_mux[26][6] , \read_value_mux[26][5] , 
        \read_value_mux[26][4] , \read_value_mux[26][3] , 
        \read_value_mux[26][2] , \read_value_mux[26][1] , 
        \read_value_mux[26][0] }) );
  cam_word_27 \words[27]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[27]), .write(write), .dec_write_index(
        dec_write_index[27]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[27]), 
        .read_results(read_results[27]), .read_value({\read_value_mux[27][31] , 
        \read_value_mux[27][30] , \read_value_mux[27][29] , 
        \read_value_mux[27][28] , \read_value_mux[27][27] , 
        \read_value_mux[27][26] , \read_value_mux[27][25] , 
        \read_value_mux[27][24] , \read_value_mux[27][23] , 
        \read_value_mux[27][22] , \read_value_mux[27][21] , 
        \read_value_mux[27][20] , \read_value_mux[27][19] , 
        \read_value_mux[27][18] , \read_value_mux[27][17] , 
        \read_value_mux[27][16] , \read_value_mux[27][15] , 
        \read_value_mux[27][14] , \read_value_mux[27][13] , 
        \read_value_mux[27][12] , \read_value_mux[27][11] , 
        \read_value_mux[27][10] , \read_value_mux[27][9] , 
        \read_value_mux[27][8] , \read_value_mux[27][7] , 
        \read_value_mux[27][6] , \read_value_mux[27][5] , 
        \read_value_mux[27][4] , \read_value_mux[27][3] , 
        \read_value_mux[27][2] , \read_value_mux[27][1] , 
        \read_value_mux[27][0] }) );
  cam_word_28 \words[28]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[28]), .write(write), .dec_write_index(
        dec_write_index[28]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[28]), 
        .read_results(read_results[28]), .read_value({\read_value_mux[28][31] , 
        \read_value_mux[28][30] , \read_value_mux[28][29] , 
        \read_value_mux[28][28] , \read_value_mux[28][27] , 
        \read_value_mux[28][26] , \read_value_mux[28][25] , 
        \read_value_mux[28][24] , \read_value_mux[28][23] , 
        \read_value_mux[28][22] , \read_value_mux[28][21] , 
        \read_value_mux[28][20] , \read_value_mux[28][19] , 
        \read_value_mux[28][18] , \read_value_mux[28][17] , 
        \read_value_mux[28][16] , \read_value_mux[28][15] , 
        \read_value_mux[28][14] , \read_value_mux[28][13] , 
        \read_value_mux[28][12] , \read_value_mux[28][11] , 
        \read_value_mux[28][10] , \read_value_mux[28][9] , 
        \read_value_mux[28][8] , \read_value_mux[28][7] , 
        \read_value_mux[28][6] , \read_value_mux[28][5] , 
        \read_value_mux[28][4] , \read_value_mux[28][3] , 
        \read_value_mux[28][2] , \read_value_mux[28][1] , 
        \read_value_mux[28][0] }) );
  cam_word_29 \words[29]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[29]), .write(write), .dec_write_index(
        dec_write_index[29]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[29]), 
        .read_results(read_results[29]), .read_value({\read_value_mux[29][31] , 
        \read_value_mux[29][30] , \read_value_mux[29][29] , 
        \read_value_mux[29][28] , \read_value_mux[29][27] , 
        \read_value_mux[29][26] , \read_value_mux[29][25] , 
        \read_value_mux[29][24] , \read_value_mux[29][23] , 
        \read_value_mux[29][22] , \read_value_mux[29][21] , 
        \read_value_mux[29][20] , \read_value_mux[29][19] , 
        \read_value_mux[29][18] , \read_value_mux[29][17] , 
        \read_value_mux[29][16] , \read_value_mux[29][15] , 
        \read_value_mux[29][14] , \read_value_mux[29][13] , 
        \read_value_mux[29][12] , \read_value_mux[29][11] , 
        \read_value_mux[29][10] , \read_value_mux[29][9] , 
        \read_value_mux[29][8] , \read_value_mux[29][7] , 
        \read_value_mux[29][6] , \read_value_mux[29][5] , 
        \read_value_mux[29][4] , \read_value_mux[29][3] , 
        \read_value_mux[29][2] , \read_value_mux[29][1] , 
        \read_value_mux[29][0] }) );
  cam_word_30 \words[30]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[30]), .write(write), .dec_write_index(
        dec_write_index[30]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[30]), 
        .read_results(read_results[30]), .read_value({\read_value_mux[30][31] , 
        \read_value_mux[30][30] , \read_value_mux[30][29] , 
        \read_value_mux[30][28] , \read_value_mux[30][27] , 
        \read_value_mux[30][26] , \read_value_mux[30][25] , 
        \read_value_mux[30][24] , \read_value_mux[30][23] , 
        \read_value_mux[30][22] , \read_value_mux[30][21] , 
        \read_value_mux[30][20] , \read_value_mux[30][19] , 
        \read_value_mux[30][18] , \read_value_mux[30][17] , 
        \read_value_mux[30][16] , \read_value_mux[30][15] , 
        \read_value_mux[30][14] , \read_value_mux[30][13] , 
        \read_value_mux[30][12] , \read_value_mux[30][11] , 
        \read_value_mux[30][10] , \read_value_mux[30][9] , 
        \read_value_mux[30][8] , \read_value_mux[30][7] , 
        \read_value_mux[30][6] , \read_value_mux[30][5] , 
        \read_value_mux[30][4] , \read_value_mux[30][3] , 
        \read_value_mux[30][2] , \read_value_mux[30][1] , 
        \read_value_mux[30][0] }) );
  cam_word_31 \words[31]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[31]), .write(write), .dec_write_index(
        dec_write_index[31]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[31]), 
        .read_results(read_results[31]), .read_value({\read_value_mux[31][31] , 
        \read_value_mux[31][30] , \read_value_mux[31][29] , 
        \read_value_mux[31][28] , \read_value_mux[31][27] , 
        \read_value_mux[31][26] , \read_value_mux[31][25] , 
        \read_value_mux[31][24] , \read_value_mux[31][23] , 
        \read_value_mux[31][22] , \read_value_mux[31][21] , 
        \read_value_mux[31][20] , \read_value_mux[31][19] , 
        \read_value_mux[31][18] , \read_value_mux[31][17] , 
        \read_value_mux[31][16] , \read_value_mux[31][15] , 
        \read_value_mux[31][14] , \read_value_mux[31][13] , 
        \read_value_mux[31][12] , \read_value_mux[31][11] , 
        \read_value_mux[31][10] , \read_value_mux[31][9] , 
        \read_value_mux[31][8] , \read_value_mux[31][7] , 
        \read_value_mux[31][6] , \read_value_mux[31][5] , 
        \read_value_mux[31][4] , \read_value_mux[31][3] , 
        \read_value_mux[31][2] , \read_value_mux[31][1] , 
        \read_value_mux[31][0] }) );
  decoder_5_32_1 read_dcdr ( .decoder_i(read_index), .decoder_o(dec_read_index) );
  decoder_5_32_0 write_dcdr ( .decoder_i(write_index), .decoder_o(
        dec_write_index) );
  priority_encoder search_ecdr ( .inp_i(search_results), .out_o(search_index), 
        .valid_o(n40) );
  mux read_mux ( .data_i({\read_value_mux[31][31] , \read_value_mux[31][30] , 
        \read_value_mux[31][29] , \read_value_mux[31][28] , 
        \read_value_mux[31][27] , \read_value_mux[31][26] , 
        \read_value_mux[31][25] , \read_value_mux[31][24] , 
        \read_value_mux[31][23] , \read_value_mux[31][22] , 
        \read_value_mux[31][21] , \read_value_mux[31][20] , 
        \read_value_mux[31][19] , \read_value_mux[31][18] , 
        \read_value_mux[31][17] , \read_value_mux[31][16] , 
        \read_value_mux[31][15] , \read_value_mux[31][14] , 
        \read_value_mux[31][13] , \read_value_mux[31][12] , 
        \read_value_mux[31][11] , \read_value_mux[31][10] , 
        \read_value_mux[31][9] , \read_value_mux[31][8] , 
        \read_value_mux[31][7] , \read_value_mux[31][6] , 
        \read_value_mux[31][5] , \read_value_mux[31][4] , 
        \read_value_mux[31][3] , \read_value_mux[31][2] , 
        \read_value_mux[31][1] , \read_value_mux[31][0] , 
        \read_value_mux[30][31] , \read_value_mux[30][30] , 
        \read_value_mux[30][29] , \read_value_mux[30][28] , 
        \read_value_mux[30][27] , \read_value_mux[30][26] , 
        \read_value_mux[30][25] , \read_value_mux[30][24] , 
        \read_value_mux[30][23] , \read_value_mux[30][22] , 
        \read_value_mux[30][21] , \read_value_mux[30][20] , 
        \read_value_mux[30][19] , \read_value_mux[30][18] , 
        \read_value_mux[30][17] , \read_value_mux[30][16] , 
        \read_value_mux[30][15] , \read_value_mux[30][14] , 
        \read_value_mux[30][13] , \read_value_mux[30][12] , 
        \read_value_mux[30][11] , \read_value_mux[30][10] , 
        \read_value_mux[30][9] , \read_value_mux[30][8] , 
        \read_value_mux[30][7] , \read_value_mux[30][6] , 
        \read_value_mux[30][5] , \read_value_mux[30][4] , 
        \read_value_mux[30][3] , \read_value_mux[30][2] , 
        \read_value_mux[30][1] , \read_value_mux[30][0] , 
        \read_value_mux[29][31] , \read_value_mux[29][30] , 
        \read_value_mux[29][29] , \read_value_mux[29][28] , 
        \read_value_mux[29][27] , \read_value_mux[29][26] , 
        \read_value_mux[29][25] , \read_value_mux[29][24] , 
        \read_value_mux[29][23] , \read_value_mux[29][22] , 
        \read_value_mux[29][21] , \read_value_mux[29][20] , 
        \read_value_mux[29][19] , \read_value_mux[29][18] , 
        \read_value_mux[29][17] , \read_value_mux[29][16] , 
        \read_value_mux[29][15] , \read_value_mux[29][14] , 
        \read_value_mux[29][13] , \read_value_mux[29][12] , 
        \read_value_mux[29][11] , \read_value_mux[29][10] , 
        \read_value_mux[29][9] , \read_value_mux[29][8] , 
        \read_value_mux[29][7] , \read_value_mux[29][6] , 
        \read_value_mux[29][5] , \read_value_mux[29][4] , 
        \read_value_mux[29][3] , \read_value_mux[29][2] , 
        \read_value_mux[29][1] , \read_value_mux[29][0] , 
        \read_value_mux[28][31] , \read_value_mux[28][30] , 
        \read_value_mux[28][29] , \read_value_mux[28][28] , 
        \read_value_mux[28][27] , \read_value_mux[28][26] , 
        \read_value_mux[28][25] , \read_value_mux[28][24] , 
        \read_value_mux[28][23] , \read_value_mux[28][22] , 
        \read_value_mux[28][21] , \read_value_mux[28][20] , 
        \read_value_mux[28][19] , \read_value_mux[28][18] , 
        \read_value_mux[28][17] , \read_value_mux[28][16] , 
        \read_value_mux[28][15] , \read_value_mux[28][14] , 
        \read_value_mux[28][13] , \read_value_mux[28][12] , 
        \read_value_mux[28][11] , \read_value_mux[28][10] , 
        \read_value_mux[28][9] , \read_value_mux[28][8] , 
        \read_value_mux[28][7] , \read_value_mux[28][6] , 
        \read_value_mux[28][5] , \read_value_mux[28][4] , 
        \read_value_mux[28][3] , \read_value_mux[28][2] , 
        \read_value_mux[28][1] , \read_value_mux[28][0] , 
        \read_value_mux[27][31] , \read_value_mux[27][30] , 
        \read_value_mux[27][29] , \read_value_mux[27][28] , 
        \read_value_mux[27][27] , \read_value_mux[27][26] , 
        \read_value_mux[27][25] , \read_value_mux[27][24] , 
        \read_value_mux[27][23] , \read_value_mux[27][22] , 
        \read_value_mux[27][21] , \read_value_mux[27][20] , 
        \read_value_mux[27][19] , \read_value_mux[27][18] , 
        \read_value_mux[27][17] , \read_value_mux[27][16] , 
        \read_value_mux[27][15] , \read_value_mux[27][14] , 
        \read_value_mux[27][13] , \read_value_mux[27][12] , 
        \read_value_mux[27][11] , \read_value_mux[27][10] , 
        \read_value_mux[27][9] , \read_value_mux[27][8] , 
        \read_value_mux[27][7] , \read_value_mux[27][6] , 
        \read_value_mux[27][5] , \read_value_mux[27][4] , 
        \read_value_mux[27][3] , \read_value_mux[27][2] , 
        \read_value_mux[27][1] , \read_value_mux[27][0] , 
        \read_value_mux[26][31] , \read_value_mux[26][30] , 
        \read_value_mux[26][29] , \read_value_mux[26][28] , 
        \read_value_mux[26][27] , \read_value_mux[26][26] , 
        \read_value_mux[26][25] , \read_value_mux[26][24] , 
        \read_value_mux[26][23] , \read_value_mux[26][22] , 
        \read_value_mux[26][21] , \read_value_mux[26][20] , 
        \read_value_mux[26][19] , \read_value_mux[26][18] , 
        \read_value_mux[26][17] , \read_value_mux[26][16] , 
        \read_value_mux[26][15] , \read_value_mux[26][14] , 
        \read_value_mux[26][13] , \read_value_mux[26][12] , 
        \read_value_mux[26][11] , \read_value_mux[26][10] , 
        \read_value_mux[26][9] , \read_value_mux[26][8] , 
        \read_value_mux[26][7] , \read_value_mux[26][6] , 
        \read_value_mux[26][5] , \read_value_mux[26][4] , 
        \read_value_mux[26][3] , \read_value_mux[26][2] , 
        \read_value_mux[26][1] , \read_value_mux[26][0] , 
        \read_value_mux[25][31] , \read_value_mux[25][30] , 
        \read_value_mux[25][29] , \read_value_mux[25][28] , 
        \read_value_mux[25][27] , \read_value_mux[25][26] , 
        \read_value_mux[25][25] , \read_value_mux[25][24] , 
        \read_value_mux[25][23] , \read_value_mux[25][22] , 
        \read_value_mux[25][21] , \read_value_mux[25][20] , 
        \read_value_mux[25][19] , \read_value_mux[25][18] , 
        \read_value_mux[25][17] , \read_value_mux[25][16] , 
        \read_value_mux[25][15] , \read_value_mux[25][14] , 
        \read_value_mux[25][13] , \read_value_mux[25][12] , 
        \read_value_mux[25][11] , \read_value_mux[25][10] , 
        \read_value_mux[25][9] , \read_value_mux[25][8] , 
        \read_value_mux[25][7] , \read_value_mux[25][6] , 
        \read_value_mux[25][5] , \read_value_mux[25][4] , 
        \read_value_mux[25][3] , \read_value_mux[25][2] , 
        \read_value_mux[25][1] , \read_value_mux[25][0] , 
        \read_value_mux[24][31] , \read_value_mux[24][30] , 
        \read_value_mux[24][29] , \read_value_mux[24][28] , 
        \read_value_mux[24][27] , \read_value_mux[24][26] , 
        \read_value_mux[24][25] , \read_value_mux[24][24] , 
        \read_value_mux[24][23] , \read_value_mux[24][22] , 
        \read_value_mux[24][21] , \read_value_mux[24][20] , 
        \read_value_mux[24][19] , \read_value_mux[24][18] , 
        \read_value_mux[24][17] , \read_value_mux[24][16] , 
        \read_value_mux[24][15] , \read_value_mux[24][14] , 
        \read_value_mux[24][13] , \read_value_mux[24][12] , 
        \read_value_mux[24][11] , \read_value_mux[24][10] , 
        \read_value_mux[24][9] , \read_value_mux[24][8] , 
        \read_value_mux[24][7] , \read_value_mux[24][6] , 
        \read_value_mux[24][5] , \read_value_mux[24][4] , 
        \read_value_mux[24][3] , \read_value_mux[24][2] , 
        \read_value_mux[24][1] , \read_value_mux[24][0] , 
        \read_value_mux[23][31] , \read_value_mux[23][30] , 
        \read_value_mux[23][29] , \read_value_mux[23][28] , 
        \read_value_mux[23][27] , \read_value_mux[23][26] , 
        \read_value_mux[23][25] , \read_value_mux[23][24] , 
        \read_value_mux[23][23] , \read_value_mux[23][22] , 
        \read_value_mux[23][21] , \read_value_mux[23][20] , 
        \read_value_mux[23][19] , \read_value_mux[23][18] , 
        \read_value_mux[23][17] , \read_value_mux[23][16] , 
        \read_value_mux[23][15] , \read_value_mux[23][14] , 
        \read_value_mux[23][13] , \read_value_mux[23][12] , 
        \read_value_mux[23][11] , \read_value_mux[23][10] , 
        \read_value_mux[23][9] , \read_value_mux[23][8] , 
        \read_value_mux[23][7] , \read_value_mux[23][6] , 
        \read_value_mux[23][5] , \read_value_mux[23][4] , 
        \read_value_mux[23][3] , \read_value_mux[23][2] , 
        \read_value_mux[23][1] , \read_value_mux[23][0] , 
        \read_value_mux[22][31] , \read_value_mux[22][30] , 
        \read_value_mux[22][29] , \read_value_mux[22][28] , 
        \read_value_mux[22][27] , \read_value_mux[22][26] , 
        \read_value_mux[22][25] , \read_value_mux[22][24] , 
        \read_value_mux[22][23] , \read_value_mux[22][22] , 
        \read_value_mux[22][21] , \read_value_mux[22][20] , 
        \read_value_mux[22][19] , \read_value_mux[22][18] , 
        \read_value_mux[22][17] , \read_value_mux[22][16] , 
        \read_value_mux[22][15] , \read_value_mux[22][14] , 
        \read_value_mux[22][13] , \read_value_mux[22][12] , 
        \read_value_mux[22][11] , \read_value_mux[22][10] , 
        \read_value_mux[22][9] , \read_value_mux[22][8] , 
        \read_value_mux[22][7] , \read_value_mux[22][6] , 
        \read_value_mux[22][5] , \read_value_mux[22][4] , 
        \read_value_mux[22][3] , \read_value_mux[22][2] , 
        \read_value_mux[22][1] , \read_value_mux[22][0] , 
        \read_value_mux[21][31] , \read_value_mux[21][30] , 
        \read_value_mux[21][29] , \read_value_mux[21][28] , 
        \read_value_mux[21][27] , \read_value_mux[21][26] , 
        \read_value_mux[21][25] , \read_value_mux[21][24] , 
        \read_value_mux[21][23] , \read_value_mux[21][22] , 
        \read_value_mux[21][21] , \read_value_mux[21][20] , 
        \read_value_mux[21][19] , \read_value_mux[21][18] , 
        \read_value_mux[21][17] , \read_value_mux[21][16] , 
        \read_value_mux[21][15] , \read_value_mux[21][14] , 
        \read_value_mux[21][13] , \read_value_mux[21][12] , 
        \read_value_mux[21][11] , \read_value_mux[21][10] , 
        \read_value_mux[21][9] , \read_value_mux[21][8] , 
        \read_value_mux[21][7] , \read_value_mux[21][6] , 
        \read_value_mux[21][5] , \read_value_mux[21][4] , 
        \read_value_mux[21][3] , \read_value_mux[21][2] , 
        \read_value_mux[21][1] , \read_value_mux[21][0] , 
        \read_value_mux[20][31] , \read_value_mux[20][30] , 
        \read_value_mux[20][29] , \read_value_mux[20][28] , 
        \read_value_mux[20][27] , \read_value_mux[20][26] , 
        \read_value_mux[20][25] , \read_value_mux[20][24] , 
        \read_value_mux[20][23] , \read_value_mux[20][22] , 
        \read_value_mux[20][21] , \read_value_mux[20][20] , 
        \read_value_mux[20][19] , \read_value_mux[20][18] , 
        \read_value_mux[20][17] , \read_value_mux[20][16] , 
        \read_value_mux[20][15] , \read_value_mux[20][14] , 
        \read_value_mux[20][13] , \read_value_mux[20][12] , 
        \read_value_mux[20][11] , \read_value_mux[20][10] , 
        \read_value_mux[20][9] , \read_value_mux[20][8] , 
        \read_value_mux[20][7] , \read_value_mux[20][6] , 
        \read_value_mux[20][5] , \read_value_mux[20][4] , 
        \read_value_mux[20][3] , \read_value_mux[20][2] , 
        \read_value_mux[20][1] , \read_value_mux[20][0] , 
        \read_value_mux[19][31] , \read_value_mux[19][30] , 
        \read_value_mux[19][29] , \read_value_mux[19][28] , 
        \read_value_mux[19][27] , \read_value_mux[19][26] , 
        \read_value_mux[19][25] , \read_value_mux[19][24] , 
        \read_value_mux[19][23] , \read_value_mux[19][22] , 
        \read_value_mux[19][21] , \read_value_mux[19][20] , 
        \read_value_mux[19][19] , \read_value_mux[19][18] , 
        \read_value_mux[19][17] , \read_value_mux[19][16] , 
        \read_value_mux[19][15] , \read_value_mux[19][14] , 
        \read_value_mux[19][13] , \read_value_mux[19][12] , 
        \read_value_mux[19][11] , \read_value_mux[19][10] , 
        \read_value_mux[19][9] , \read_value_mux[19][8] , 
        \read_value_mux[19][7] , \read_value_mux[19][6] , 
        \read_value_mux[19][5] , \read_value_mux[19][4] , 
        \read_value_mux[19][3] , \read_value_mux[19][2] , 
        \read_value_mux[19][1] , \read_value_mux[19][0] , 
        \read_value_mux[18][31] , \read_value_mux[18][30] , 
        \read_value_mux[18][29] , \read_value_mux[18][28] , 
        \read_value_mux[18][27] , \read_value_mux[18][26] , 
        \read_value_mux[18][25] , \read_value_mux[18][24] , 
        \read_value_mux[18][23] , \read_value_mux[18][22] , 
        \read_value_mux[18][21] , \read_value_mux[18][20] , 
        \read_value_mux[18][19] , \read_value_mux[18][18] , 
        \read_value_mux[18][17] , \read_value_mux[18][16] , 
        \read_value_mux[18][15] , \read_value_mux[18][14] , 
        \read_value_mux[18][13] , \read_value_mux[18][12] , 
        \read_value_mux[18][11] , \read_value_mux[18][10] , 
        \read_value_mux[18][9] , \read_value_mux[18][8] , 
        \read_value_mux[18][7] , \read_value_mux[18][6] , 
        \read_value_mux[18][5] , \read_value_mux[18][4] , 
        \read_value_mux[18][3] , \read_value_mux[18][2] , 
        \read_value_mux[18][1] , \read_value_mux[18][0] , 
        \read_value_mux[17][31] , \read_value_mux[17][30] , 
        \read_value_mux[17][29] , \read_value_mux[17][28] , 
        \read_value_mux[17][27] , \read_value_mux[17][26] , 
        \read_value_mux[17][25] , \read_value_mux[17][24] , 
        \read_value_mux[17][23] , \read_value_mux[17][22] , 
        \read_value_mux[17][21] , \read_value_mux[17][20] , 
        \read_value_mux[17][19] , \read_value_mux[17][18] , 
        \read_value_mux[17][17] , \read_value_mux[17][16] , 
        \read_value_mux[17][15] , \read_value_mux[17][14] , 
        \read_value_mux[17][13] , \read_value_mux[17][12] , 
        \read_value_mux[17][11] , \read_value_mux[17][10] , 
        \read_value_mux[17][9] , \read_value_mux[17][8] , 
        \read_value_mux[17][7] , \read_value_mux[17][6] , 
        \read_value_mux[17][5] , \read_value_mux[17][4] , 
        \read_value_mux[17][3] , \read_value_mux[17][2] , 
        \read_value_mux[17][1] , \read_value_mux[17][0] , 
        \read_value_mux[16][31] , \read_value_mux[16][30] , 
        \read_value_mux[16][29] , \read_value_mux[16][28] , 
        \read_value_mux[16][27] , \read_value_mux[16][26] , 
        \read_value_mux[16][25] , \read_value_mux[16][24] , 
        \read_value_mux[16][23] , \read_value_mux[16][22] , 
        \read_value_mux[16][21] , \read_value_mux[16][20] , 
        \read_value_mux[16][19] , \read_value_mux[16][18] , 
        \read_value_mux[16][17] , \read_value_mux[16][16] , 
        \read_value_mux[16][15] , \read_value_mux[16][14] , 
        \read_value_mux[16][13] , \read_value_mux[16][12] , 
        \read_value_mux[16][11] , \read_value_mux[16][10] , 
        \read_value_mux[16][9] , \read_value_mux[16][8] , 
        \read_value_mux[16][7] , \read_value_mux[16][6] , 
        \read_value_mux[16][5] , \read_value_mux[16][4] , 
        \read_value_mux[16][3] , \read_value_mux[16][2] , 
        \read_value_mux[16][1] , \read_value_mux[16][0] , 
        \read_value_mux[15][31] , \read_value_mux[15][30] , 
        \read_value_mux[15][29] , \read_value_mux[15][28] , 
        \read_value_mux[15][27] , \read_value_mux[15][26] , 
        \read_value_mux[15][25] , \read_value_mux[15][24] , 
        \read_value_mux[15][23] , \read_value_mux[15][22] , 
        \read_value_mux[15][21] , \read_value_mux[15][20] , 
        \read_value_mux[15][19] , \read_value_mux[15][18] , 
        \read_value_mux[15][17] , \read_value_mux[15][16] , 
        \read_value_mux[15][15] , \read_value_mux[15][14] , 
        \read_value_mux[15][13] , \read_value_mux[15][12] , 
        \read_value_mux[15][11] , \read_value_mux[15][10] , 
        \read_value_mux[15][9] , \read_value_mux[15][8] , 
        \read_value_mux[15][7] , \read_value_mux[15][6] , 
        \read_value_mux[15][5] , \read_value_mux[15][4] , 
        \read_value_mux[15][3] , \read_value_mux[15][2] , 
        \read_value_mux[15][1] , \read_value_mux[15][0] , 
        \read_value_mux[14][31] , \read_value_mux[14][30] , 
        \read_value_mux[14][29] , \read_value_mux[14][28] , 
        \read_value_mux[14][27] , \read_value_mux[14][26] , 
        \read_value_mux[14][25] , \read_value_mux[14][24] , 
        \read_value_mux[14][23] , \read_value_mux[14][22] , 
        \read_value_mux[14][21] , \read_value_mux[14][20] , 
        \read_value_mux[14][19] , \read_value_mux[14][18] , 
        \read_value_mux[14][17] , \read_value_mux[14][16] , 
        \read_value_mux[14][15] , \read_value_mux[14][14] , 
        \read_value_mux[14][13] , \read_value_mux[14][12] , 
        \read_value_mux[14][11] , \read_value_mux[14][10] , 
        \read_value_mux[14][9] , \read_value_mux[14][8] , 
        \read_value_mux[14][7] , \read_value_mux[14][6] , 
        \read_value_mux[14][5] , \read_value_mux[14][4] , 
        \read_value_mux[14][3] , \read_value_mux[14][2] , 
        \read_value_mux[14][1] , \read_value_mux[14][0] , 
        \read_value_mux[13][31] , \read_value_mux[13][30] , 
        \read_value_mux[13][29] , \read_value_mux[13][28] , 
        \read_value_mux[13][27] , \read_value_mux[13][26] , 
        \read_value_mux[13][25] , \read_value_mux[13][24] , 
        \read_value_mux[13][23] , \read_value_mux[13][22] , 
        \read_value_mux[13][21] , \read_value_mux[13][20] , 
        \read_value_mux[13][19] , \read_value_mux[13][18] , 
        \read_value_mux[13][17] , \read_value_mux[13][16] , 
        \read_value_mux[13][15] , \read_value_mux[13][14] , 
        \read_value_mux[13][13] , \read_value_mux[13][12] , 
        \read_value_mux[13][11] , \read_value_mux[13][10] , 
        \read_value_mux[13][9] , \read_value_mux[13][8] , 
        \read_value_mux[13][7] , \read_value_mux[13][6] , 
        \read_value_mux[13][5] , \read_value_mux[13][4] , 
        \read_value_mux[13][3] , \read_value_mux[13][2] , 
        \read_value_mux[13][1] , \read_value_mux[13][0] , 
        \read_value_mux[12][31] , \read_value_mux[12][30] , 
        \read_value_mux[12][29] , \read_value_mux[12][28] , 
        \read_value_mux[12][27] , \read_value_mux[12][26] , 
        \read_value_mux[12][25] , \read_value_mux[12][24] , 
        \read_value_mux[12][23] , \read_value_mux[12][22] , 
        \read_value_mux[12][21] , \read_value_mux[12][20] , 
        \read_value_mux[12][19] , \read_value_mux[12][18] , 
        \read_value_mux[12][17] , \read_value_mux[12][16] , 
        \read_value_mux[12][15] , \read_value_mux[12][14] , 
        \read_value_mux[12][13] , \read_value_mux[12][12] , 
        \read_value_mux[12][11] , \read_value_mux[12][10] , 
        \read_value_mux[12][9] , \read_value_mux[12][8] , 
        \read_value_mux[12][7] , \read_value_mux[12][6] , 
        \read_value_mux[12][5] , \read_value_mux[12][4] , 
        \read_value_mux[12][3] , \read_value_mux[12][2] , 
        \read_value_mux[12][1] , \read_value_mux[12][0] , 
        \read_value_mux[11][31] , \read_value_mux[11][30] , 
        \read_value_mux[11][29] , \read_value_mux[11][28] , 
        \read_value_mux[11][27] , \read_value_mux[11][26] , 
        \read_value_mux[11][25] , \read_value_mux[11][24] , 
        \read_value_mux[11][23] , \read_value_mux[11][22] , 
        \read_value_mux[11][21] , \read_value_mux[11][20] , 
        \read_value_mux[11][19] , \read_value_mux[11][18] , 
        \read_value_mux[11][17] , \read_value_mux[11][16] , 
        \read_value_mux[11][15] , \read_value_mux[11][14] , 
        \read_value_mux[11][13] , \read_value_mux[11][12] , 
        \read_value_mux[11][11] , \read_value_mux[11][10] , 
        \read_value_mux[11][9] , \read_value_mux[11][8] , 
        \read_value_mux[11][7] , \read_value_mux[11][6] , 
        \read_value_mux[11][5] , \read_value_mux[11][4] , 
        \read_value_mux[11][3] , \read_value_mux[11][2] , 
        \read_value_mux[11][1] , \read_value_mux[11][0] , 
        \read_value_mux[10][31] , \read_value_mux[10][30] , 
        \read_value_mux[10][29] , \read_value_mux[10][28] , 
        \read_value_mux[10][27] , \read_value_mux[10][26] , 
        \read_value_mux[10][25] , \read_value_mux[10][24] , 
        \read_value_mux[10][23] , \read_value_mux[10][22] , 
        \read_value_mux[10][21] , \read_value_mux[10][20] , 
        \read_value_mux[10][19] , \read_value_mux[10][18] , 
        \read_value_mux[10][17] , \read_value_mux[10][16] , 
        \read_value_mux[10][15] , \read_value_mux[10][14] , 
        \read_value_mux[10][13] , \read_value_mux[10][12] , 
        \read_value_mux[10][11] , \read_value_mux[10][10] , 
        \read_value_mux[10][9] , \read_value_mux[10][8] , 
        \read_value_mux[10][7] , \read_value_mux[10][6] , 
        \read_value_mux[10][5] , \read_value_mux[10][4] , 
        \read_value_mux[10][3] , \read_value_mux[10][2] , 
        \read_value_mux[10][1] , \read_value_mux[10][0] , 
        \read_value_mux[9][31] , \read_value_mux[9][30] , 
        \read_value_mux[9][29] , \read_value_mux[9][28] , 
        \read_value_mux[9][27] , \read_value_mux[9][26] , 
        \read_value_mux[9][25] , \read_value_mux[9][24] , 
        \read_value_mux[9][23] , \read_value_mux[9][22] , 
        \read_value_mux[9][21] , \read_value_mux[9][20] , 
        \read_value_mux[9][19] , \read_value_mux[9][18] , 
        \read_value_mux[9][17] , \read_value_mux[9][16] , 
        \read_value_mux[9][15] , \read_value_mux[9][14] , 
        \read_value_mux[9][13] , \read_value_mux[9][12] , 
        \read_value_mux[9][11] , \read_value_mux[9][10] , 
        \read_value_mux[9][9] , \read_value_mux[9][8] , \read_value_mux[9][7] , 
        \read_value_mux[9][6] , \read_value_mux[9][5] , \read_value_mux[9][4] , 
        \read_value_mux[9][3] , \read_value_mux[9][2] , \read_value_mux[9][1] , 
        \read_value_mux[9][0] , \read_value_mux[8][31] , 
        \read_value_mux[8][30] , \read_value_mux[8][29] , 
        \read_value_mux[8][28] , \read_value_mux[8][27] , 
        \read_value_mux[8][26] , \read_value_mux[8][25] , 
        \read_value_mux[8][24] , \read_value_mux[8][23] , 
        \read_value_mux[8][22] , \read_value_mux[8][21] , 
        \read_value_mux[8][20] , \read_value_mux[8][19] , 
        \read_value_mux[8][18] , \read_value_mux[8][17] , 
        \read_value_mux[8][16] , \read_value_mux[8][15] , 
        \read_value_mux[8][14] , \read_value_mux[8][13] , 
        \read_value_mux[8][12] , \read_value_mux[8][11] , 
        \read_value_mux[8][10] , \read_value_mux[8][9] , 
        \read_value_mux[8][8] , \read_value_mux[8][7] , \read_value_mux[8][6] , 
        \read_value_mux[8][5] , \read_value_mux[8][4] , \read_value_mux[8][3] , 
        \read_value_mux[8][2] , \read_value_mux[8][1] , \read_value_mux[8][0] , 
        \read_value_mux[7][31] , \read_value_mux[7][30] , 
        \read_value_mux[7][29] , \read_value_mux[7][28] , 
        \read_value_mux[7][27] , \read_value_mux[7][26] , 
        \read_value_mux[7][25] , \read_value_mux[7][24] , 
        \read_value_mux[7][23] , \read_value_mux[7][22] , 
        \read_value_mux[7][21] , \read_value_mux[7][20] , 
        \read_value_mux[7][19] , \read_value_mux[7][18] , 
        \read_value_mux[7][17] , \read_value_mux[7][16] , 
        \read_value_mux[7][15] , \read_value_mux[7][14] , 
        \read_value_mux[7][13] , \read_value_mux[7][12] , 
        \read_value_mux[7][11] , \read_value_mux[7][10] , 
        \read_value_mux[7][9] , \read_value_mux[7][8] , \read_value_mux[7][7] , 
        \read_value_mux[7][6] , \read_value_mux[7][5] , \read_value_mux[7][4] , 
        \read_value_mux[7][3] , \read_value_mux[7][2] , \read_value_mux[7][1] , 
        \read_value_mux[7][0] , \read_value_mux[6][31] , 
        \read_value_mux[6][30] , \read_value_mux[6][29] , 
        \read_value_mux[6][28] , \read_value_mux[6][27] , 
        \read_value_mux[6][26] , \read_value_mux[6][25] , 
        \read_value_mux[6][24] , \read_value_mux[6][23] , 
        \read_value_mux[6][22] , \read_value_mux[6][21] , 
        \read_value_mux[6][20] , \read_value_mux[6][19] , 
        \read_value_mux[6][18] , \read_value_mux[6][17] , 
        \read_value_mux[6][16] , \read_value_mux[6][15] , 
        \read_value_mux[6][14] , \read_value_mux[6][13] , 
        \read_value_mux[6][12] , \read_value_mux[6][11] , 
        \read_value_mux[6][10] , \read_value_mux[6][9] , 
        \read_value_mux[6][8] , \read_value_mux[6][7] , \read_value_mux[6][6] , 
        \read_value_mux[6][5] , \read_value_mux[6][4] , \read_value_mux[6][3] , 
        \read_value_mux[6][2] , \read_value_mux[6][1] , \read_value_mux[6][0] , 
        \read_value_mux[5][31] , \read_value_mux[5][30] , 
        \read_value_mux[5][29] , \read_value_mux[5][28] , 
        \read_value_mux[5][27] , \read_value_mux[5][26] , 
        \read_value_mux[5][25] , \read_value_mux[5][24] , 
        \read_value_mux[5][23] , \read_value_mux[5][22] , 
        \read_value_mux[5][21] , \read_value_mux[5][20] , 
        \read_value_mux[5][19] , \read_value_mux[5][18] , 
        \read_value_mux[5][17] , \read_value_mux[5][16] , 
        \read_value_mux[5][15] , \read_value_mux[5][14] , 
        \read_value_mux[5][13] , \read_value_mux[5][12] , 
        \read_value_mux[5][11] , \read_value_mux[5][10] , 
        \read_value_mux[5][9] , \read_value_mux[5][8] , \read_value_mux[5][7] , 
        \read_value_mux[5][6] , \read_value_mux[5][5] , \read_value_mux[5][4] , 
        \read_value_mux[5][3] , \read_value_mux[5][2] , \read_value_mux[5][1] , 
        \read_value_mux[5][0] , \read_value_mux[4][31] , 
        \read_value_mux[4][30] , \read_value_mux[4][29] , 
        \read_value_mux[4][28] , \read_value_mux[4][27] , 
        \read_value_mux[4][26] , \read_value_mux[4][25] , 
        \read_value_mux[4][24] , \read_value_mux[4][23] , 
        \read_value_mux[4][22] , \read_value_mux[4][21] , 
        \read_value_mux[4][20] , \read_value_mux[4][19] , 
        \read_value_mux[4][18] , \read_value_mux[4][17] , 
        \read_value_mux[4][16] , \read_value_mux[4][15] , 
        \read_value_mux[4][14] , \read_value_mux[4][13] , 
        \read_value_mux[4][12] , \read_value_mux[4][11] , 
        \read_value_mux[4][10] , \read_value_mux[4][9] , 
        \read_value_mux[4][8] , \read_value_mux[4][7] , \read_value_mux[4][6] , 
        \read_value_mux[4][5] , \read_value_mux[4][4] , \read_value_mux[4][3] , 
        \read_value_mux[4][2] , \read_value_mux[4][1] , \read_value_mux[4][0] , 
        \read_value_mux[3][31] , \read_value_mux[3][30] , 
        \read_value_mux[3][29] , \read_value_mux[3][28] , 
        \read_value_mux[3][27] , \read_value_mux[3][26] , 
        \read_value_mux[3][25] , \read_value_mux[3][24] , 
        \read_value_mux[3][23] , \read_value_mux[3][22] , 
        \read_value_mux[3][21] , \read_value_mux[3][20] , 
        \read_value_mux[3][19] , \read_value_mux[3][18] , 
        \read_value_mux[3][17] , \read_value_mux[3][16] , 
        \read_value_mux[3][15] , \read_value_mux[3][14] , 
        \read_value_mux[3][13] , \read_value_mux[3][12] , 
        \read_value_mux[3][11] , \read_value_mux[3][10] , 
        \read_value_mux[3][9] , \read_value_mux[3][8] , \read_value_mux[3][7] , 
        \read_value_mux[3][6] , \read_value_mux[3][5] , \read_value_mux[3][4] , 
        \read_value_mux[3][3] , \read_value_mux[3][2] , \read_value_mux[3][1] , 
        \read_value_mux[3][0] , \read_value_mux[2][31] , 
        \read_value_mux[2][30] , \read_value_mux[2][29] , 
        \read_value_mux[2][28] , \read_value_mux[2][27] , 
        \read_value_mux[2][26] , \read_value_mux[2][25] , 
        \read_value_mux[2][24] , \read_value_mux[2][23] , 
        \read_value_mux[2][22] , \read_value_mux[2][21] , 
        \read_value_mux[2][20] , \read_value_mux[2][19] , 
        \read_value_mux[2][18] , \read_value_mux[2][17] , 
        \read_value_mux[2][16] , \read_value_mux[2][15] , 
        \read_value_mux[2][14] , \read_value_mux[2][13] , 
        \read_value_mux[2][12] , \read_value_mux[2][11] , 
        \read_value_mux[2][10] , \read_value_mux[2][9] , 
        \read_value_mux[2][8] , \read_value_mux[2][7] , \read_value_mux[2][6] , 
        \read_value_mux[2][5] , \read_value_mux[2][4] , \read_value_mux[2][3] , 
        \read_value_mux[2][2] , \read_value_mux[2][1] , \read_value_mux[2][0] , 
        \read_value_mux[1][31] , \read_value_mux[1][30] , 
        \read_value_mux[1][29] , \read_value_mux[1][28] , 
        \read_value_mux[1][27] , \read_value_mux[1][26] , 
        \read_value_mux[1][25] , \read_value_mux[1][24] , 
        \read_value_mux[1][23] , \read_value_mux[1][22] , 
        \read_value_mux[1][21] , \read_value_mux[1][20] , 
        \read_value_mux[1][19] , \read_value_mux[1][18] , 
        \read_value_mux[1][17] , \read_value_mux[1][16] , 
        \read_value_mux[1][15] , \read_value_mux[1][14] , 
        \read_value_mux[1][13] , \read_value_mux[1][12] , 
        \read_value_mux[1][11] , \read_value_mux[1][10] , 
        \read_value_mux[1][9] , \read_value_mux[1][8] , \read_value_mux[1][7] , 
        \read_value_mux[1][6] , \read_value_mux[1][5] , \read_value_mux[1][4] , 
        \read_value_mux[1][3] , \read_value_mux[1][2] , \read_value_mux[1][1] , 
        \read_value_mux[1][0] , \read_value_mux[0][31] , 
        \read_value_mux[0][30] , \read_value_mux[0][29] , 
        \read_value_mux[0][28] , \read_value_mux[0][27] , 
        \read_value_mux[0][26] , \read_value_mux[0][25] , 
        \read_value_mux[0][24] , \read_value_mux[0][23] , 
        \read_value_mux[0][22] , \read_value_mux[0][21] , 
        \read_value_mux[0][20] , \read_value_mux[0][19] , 
        \read_value_mux[0][18] , \read_value_mux[0][17] , 
        \read_value_mux[0][16] , \read_value_mux[0][15] , 
        \read_value_mux[0][14] , \read_value_mux[0][13] , 
        \read_value_mux[0][12] , \read_value_mux[0][11] , 
        \read_value_mux[0][10] , \read_value_mux[0][9] , 
        \read_value_mux[0][8] , \read_value_mux[0][7] , \read_value_mux[0][6] , 
        \read_value_mux[0][5] , \read_value_mux[0][4] , \read_value_mux[0][3] , 
        \read_value_mux[0][2] , \read_value_mux[0][1] , \read_value_mux[0][0] }), .select_i(read_index), .data_o(read_value) );
  NR4D0 U23 ( .A1(search_results[10]), .A2(search_results[11]), .A3(
        search_results[13]), .A4(search_results[12]), .ZN(n20) );
  NR4D0 U24 ( .A1(search_results[7]), .A2(search_results[22]), .A3(
        search_results[9]), .A4(search_results[8]), .ZN(n21) );
  NR4D0 U25 ( .A1(search_results[6]), .A2(search_results[4]), .A3(
        search_results[5]), .A4(search_results[3]), .ZN(n22) );
  NR4D0 U26 ( .A1(search_results[1]), .A2(search_results[14]), .A3(
        search_results[30]), .A4(search_results[2]), .ZN(n23) );
  ND4D0 U27 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .ZN(n24) );
  NR4D0 U28 ( .A1(search_results[27]), .A2(search_results[31]), .A3(
        search_results[28]), .A4(search_results[26]), .ZN(n25) );
  NR4D0 U29 ( .A1(search_results[24]), .A2(search_results[23]), .A3(
        search_results[25]), .A4(search_results[0]), .ZN(n26) );
  NR4D0 U30 ( .A1(search_results[21]), .A2(search_results[20]), .A3(
        search_results[19]), .A4(search_results[18]), .ZN(n27) );
  NR4D0 U31 ( .A1(search_results[16]), .A2(search_results[15]), .A3(
        search_results[29]), .A4(search_results[17]), .ZN(n28) );
  ND4D0 U32 ( .A1(n25), .A2(n26), .A3(n27), .A4(n28), .ZN(n29) );
  OA21D0 U33 ( .A1(n24), .A2(n29), .B(n40), .Z(search_valid) );
  NR4D0 U34 ( .A1(read_results[31]), .A2(read_results[30]), .A3(
        read_results[29]), .A4(read_results[28]), .ZN(n30) );
  NR4D0 U35 ( .A1(read_results[27]), .A2(read_results[26]), .A3(
        read_results[25]), .A4(read_results[24]), .ZN(n31) );
  NR4D0 U36 ( .A1(read_results[23]), .A2(read_results[22]), .A3(
        read_results[21]), .A4(read_results[20]), .ZN(n32) );
  NR4D0 U37 ( .A1(read_results[19]), .A2(read_results[18]), .A3(
        read_results[17]), .A4(read_results[16]), .ZN(n33) );
  AN4D0 U38 ( .A1(n30), .A2(n31), .A3(n32), .A4(n33), .Z(n34) );
  NR4D0 U39 ( .A1(read_results[15]), .A2(read_results[14]), .A3(
        read_results[13]), .A4(read_results[12]), .ZN(n35) );
  NR4D0 U40 ( .A1(read_results[11]), .A2(read_results[10]), .A3(
        read_results[9]), .A4(read_results[8]), .ZN(n36) );
  NR4D0 U41 ( .A1(read_results[7]), .A2(read_results[6]), .A3(read_results[5]), 
        .A4(read_results[4]), .ZN(n37) );
  NR4D0 U42 ( .A1(read_results[3]), .A2(read_results[2]), .A3(read_results[1]), 
        .A4(read_results[0]), .ZN(n38) );
  AN4D0 U43 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .Z(n39) );
  CKND2D0 U44 ( .A1(n34), .A2(n39), .ZN(read_valid) );
endmodule

