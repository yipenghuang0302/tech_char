
module decoder_5_32_1 ( decoder_i, decoder_o );
  input [4:0] decoder_i;
  output [31:0] decoder_o;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96;

  GTECH_AND2 C4 ( .A(decoder_i[4]), .B(decoder_i[3]), .Z(N0) );
  GTECH_AND2 C5 ( .A(decoder_i[2]), .B(decoder_i[1]), .Z(N1) );
  GTECH_AND2 C6 ( .A(N0), .B(N1), .Z(N2) );
  GTECH_AND2 C7 ( .A(N2), .B(decoder_i[0]), .Z(N3) );
  GTECH_OR2 C17 ( .A(N88), .B(N89), .Z(N4) );
  GTECH_OR2 C18 ( .A(N90), .B(N91), .Z(N5) );
  GTECH_OR2 C19 ( .A(N4), .B(N5), .Z(N6) );
  GTECH_OR2 C20 ( .A(N6), .B(decoder_i[0]), .Z(N7) );
  GTECH_OR2 C32 ( .A(N90), .B(decoder_i[1]), .Z(N9) );
  GTECH_OR2 C33 ( .A(N4), .B(N9), .Z(N10) );
  GTECH_OR2 C34 ( .A(N10), .B(N92), .Z(N11) );
  GTECH_OR2 C47 ( .A(N10), .B(decoder_i[0]), .Z(N13) );
  GTECH_OR2 C59 ( .A(decoder_i[2]), .B(N91), .Z(N15) );
  GTECH_OR2 C60 ( .A(N4), .B(N15), .Z(N16) );
  GTECH_OR2 C61 ( .A(N16), .B(N92), .Z(N17) );
  GTECH_OR2 C74 ( .A(N16), .B(decoder_i[0]), .Z(N19) );
  GTECH_OR2 C85 ( .A(decoder_i[2]), .B(decoder_i[1]), .Z(N21) );
  GTECH_OR2 C86 ( .A(N4), .B(N21), .Z(N22) );
  GTECH_OR2 C87 ( .A(N22), .B(N92), .Z(N23) );
  GTECH_OR2 C99 ( .A(N22), .B(decoder_i[0]), .Z(N25) );
  GTECH_OR2 C110 ( .A(N88), .B(decoder_i[3]), .Z(N27) );
  GTECH_OR2 C112 ( .A(N27), .B(N5), .Z(N28) );
  GTECH_OR2 C113 ( .A(N28), .B(N92), .Z(N29) );
  GTECH_OR2 C126 ( .A(N28), .B(decoder_i[0]), .Z(N31) );
  GTECH_OR2 C138 ( .A(N27), .B(N9), .Z(N33) );
  GTECH_OR2 C139 ( .A(N33), .B(N92), .Z(N34) );
  GTECH_OR2 C151 ( .A(N33), .B(decoder_i[0]), .Z(N36) );
  GTECH_OR2 C163 ( .A(N27), .B(N15), .Z(N38) );
  GTECH_OR2 C164 ( .A(N38), .B(N92), .Z(N39) );
  GTECH_OR2 C176 ( .A(N38), .B(decoder_i[0]), .Z(N41) );
  GTECH_OR2 C187 ( .A(N27), .B(N21), .Z(N43) );
  GTECH_OR2 C188 ( .A(N43), .B(N92), .Z(N44) );
  GTECH_OR2 C199 ( .A(N43), .B(decoder_i[0]), .Z(N46) );
  GTECH_OR2 C210 ( .A(decoder_i[4]), .B(N89), .Z(N48) );
  GTECH_OR2 C212 ( .A(N48), .B(N5), .Z(N49) );
  GTECH_OR2 C213 ( .A(N49), .B(N92), .Z(N50) );
  GTECH_OR2 C226 ( .A(N49), .B(decoder_i[0]), .Z(N52) );
  GTECH_OR2 C238 ( .A(N48), .B(N9), .Z(N54) );
  GTECH_OR2 C239 ( .A(N54), .B(N92), .Z(N55) );
  GTECH_OR2 C251 ( .A(N54), .B(decoder_i[0]), .Z(N57) );
  GTECH_OR2 C263 ( .A(N48), .B(N15), .Z(N59) );
  GTECH_OR2 C264 ( .A(N59), .B(N92), .Z(N60) );
  GTECH_OR2 C276 ( .A(N59), .B(decoder_i[0]), .Z(N62) );
  GTECH_OR2 C287 ( .A(N48), .B(N21), .Z(N64) );
  GTECH_OR2 C288 ( .A(N64), .B(N92), .Z(N65) );
  GTECH_OR2 C299 ( .A(N64), .B(decoder_i[0]), .Z(N67) );
  GTECH_OR2 C309 ( .A(decoder_i[4]), .B(decoder_i[3]), .Z(N69) );
  GTECH_OR2 C311 ( .A(N69), .B(N5), .Z(N70) );
  GTECH_OR2 C312 ( .A(N70), .B(N92), .Z(N71) );
  GTECH_OR2 C324 ( .A(N70), .B(decoder_i[0]), .Z(N73) );
  GTECH_OR2 C335 ( .A(N69), .B(N9), .Z(N75) );
  GTECH_OR2 C336 ( .A(N75), .B(N92), .Z(N76) );
  GTECH_OR2 C347 ( .A(N75), .B(decoder_i[0]), .Z(N78) );
  GTECH_OR2 C358 ( .A(N69), .B(N15), .Z(N80) );
  GTECH_OR2 C359 ( .A(N80), .B(N92), .Z(N81) );
  GTECH_OR2 C370 ( .A(N80), .B(decoder_i[0]), .Z(N83) );
  GTECH_OR2 C380 ( .A(N69), .B(N21), .Z(N85) );
  GTECH_OR2 C381 ( .A(N85), .B(N92), .Z(N86) );
  GTECH_AND2 C393 ( .A(N88), .B(N89), .Z(N93) );
  GTECH_AND2 C394 ( .A(N90), .B(N91), .Z(N94) );
  GTECH_AND2 C395 ( .A(N93), .B(N94), .Z(N95) );
  GTECH_AND2 C396 ( .A(N95), .B(N92), .Z(N96) );
  GTECH_BUF B_0 ( .A(N3), .Z(decoder_o[31]) );
  GTECH_NOT I_0 ( .A(N7), .Z(N8) );
  GTECH_BUF B_1 ( .A(N8), .Z(decoder_o[30]) );
  GTECH_NOT I_1 ( .A(N11), .Z(N12) );
  GTECH_BUF B_2 ( .A(N12), .Z(decoder_o[29]) );
  GTECH_NOT I_2 ( .A(N13), .Z(N14) );
  GTECH_BUF B_3 ( .A(N14), .Z(decoder_o[28]) );
  GTECH_NOT I_3 ( .A(N17), .Z(N18) );
  GTECH_BUF B_4 ( .A(N18), .Z(decoder_o[27]) );
  GTECH_NOT I_4 ( .A(N19), .Z(N20) );
  GTECH_BUF B_5 ( .A(N20), .Z(decoder_o[26]) );
  GTECH_NOT I_5 ( .A(N23), .Z(N24) );
  GTECH_BUF B_6 ( .A(N24), .Z(decoder_o[25]) );
  GTECH_NOT I_6 ( .A(N25), .Z(N26) );
  GTECH_BUF B_7 ( .A(N26), .Z(decoder_o[24]) );
  GTECH_NOT I_7 ( .A(N29), .Z(N30) );
  GTECH_BUF B_8 ( .A(N30), .Z(decoder_o[23]) );
  GTECH_NOT I_8 ( .A(N31), .Z(N32) );
  GTECH_BUF B_9 ( .A(N32), .Z(decoder_o[22]) );
  GTECH_NOT I_9 ( .A(N34), .Z(N35) );
  GTECH_BUF B_10 ( .A(N35), .Z(decoder_o[21]) );
  GTECH_NOT I_10 ( .A(N36), .Z(N37) );
  GTECH_BUF B_11 ( .A(N37), .Z(decoder_o[20]) );
  GTECH_NOT I_11 ( .A(N39), .Z(N40) );
  GTECH_BUF B_12 ( .A(N40), .Z(decoder_o[19]) );
  GTECH_NOT I_12 ( .A(N41), .Z(N42) );
  GTECH_BUF B_13 ( .A(N42), .Z(decoder_o[18]) );
  GTECH_NOT I_13 ( .A(N44), .Z(N45) );
  GTECH_BUF B_14 ( .A(N45), .Z(decoder_o[17]) );
  GTECH_NOT I_14 ( .A(N46), .Z(N47) );
  GTECH_BUF B_15 ( .A(N47), .Z(decoder_o[16]) );
  GTECH_NOT I_15 ( .A(N50), .Z(N51) );
  GTECH_BUF B_16 ( .A(N51), .Z(decoder_o[15]) );
  GTECH_NOT I_16 ( .A(N52), .Z(N53) );
  GTECH_BUF B_17 ( .A(N53), .Z(decoder_o[14]) );
  GTECH_NOT I_17 ( .A(N55), .Z(N56) );
  GTECH_BUF B_18 ( .A(N56), .Z(decoder_o[13]) );
  GTECH_NOT I_18 ( .A(N57), .Z(N58) );
  GTECH_BUF B_19 ( .A(N58), .Z(decoder_o[12]) );
  GTECH_NOT I_19 ( .A(N60), .Z(N61) );
  GTECH_BUF B_20 ( .A(N61), .Z(decoder_o[11]) );
  GTECH_NOT I_20 ( .A(N62), .Z(N63) );
  GTECH_BUF B_21 ( .A(N63), .Z(decoder_o[10]) );
  GTECH_NOT I_21 ( .A(N65), .Z(N66) );
  GTECH_BUF B_22 ( .A(N66), .Z(decoder_o[9]) );
  GTECH_NOT I_22 ( .A(N67), .Z(N68) );
  GTECH_BUF B_23 ( .A(N68), .Z(decoder_o[8]) );
  GTECH_NOT I_23 ( .A(N71), .Z(N72) );
  GTECH_BUF B_24 ( .A(N72), .Z(decoder_o[7]) );
  GTECH_NOT I_24 ( .A(N73), .Z(N74) );
  GTECH_BUF B_25 ( .A(N74), .Z(decoder_o[6]) );
  GTECH_NOT I_25 ( .A(N76), .Z(N77) );
  GTECH_BUF B_26 ( .A(N77), .Z(decoder_o[5]) );
  GTECH_NOT I_26 ( .A(N78), .Z(N79) );
  GTECH_BUF B_27 ( .A(N79), .Z(decoder_o[4]) );
  GTECH_NOT I_27 ( .A(N81), .Z(N82) );
  GTECH_BUF B_28 ( .A(N82), .Z(decoder_o[3]) );
  GTECH_NOT I_28 ( .A(N83), .Z(N84) );
  GTECH_BUF B_29 ( .A(N84), .Z(decoder_o[2]) );
  GTECH_NOT I_29 ( .A(N86), .Z(N87) );
  GTECH_BUF B_30 ( .A(N87), .Z(decoder_o[1]) );
  GTECH_NOT I_30 ( .A(decoder_i[4]), .Z(N88) );
  GTECH_NOT I_31 ( .A(decoder_i[3]), .Z(N89) );
  GTECH_NOT I_32 ( .A(decoder_i[2]), .Z(N90) );
  GTECH_NOT I_33 ( .A(decoder_i[1]), .Z(N91) );
  GTECH_NOT I_34 ( .A(decoder_i[0]), .Z(N92) );
  GTECH_BUF B_31 ( .A(N96), .Z(decoder_o[0]) );
endmodule


module priority_encoder ( inp_i, out_o, valid_o );
  input [31:0] inp_i;
  output [4:0] out_o;
  output valid_o;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242,
         N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253,
         N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264,
         N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374,
         N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385,
         N386, N387, N388, N389, N390, N391, N392, N393, N394, N395, N396,
         N397, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440,
         N441, N442, N443, N444, N445, N446, N447, N448, N449, N450, N451,
         N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, N462,
         N463, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N496, N497, N498, N499, N500, N501, N502, N503, N504, N505, N506,
         N507, N508, N509, N510, N511, N512, N513, N514, N515, N516, N517,
         N518, N519, N520, N521, N522, N523, N524, N525, N526, N527, N528,
         N529, N530, N531, N532, N533, N534, N535, N536, N537, N538;

  GTECH_AND2 C20 ( .A(inp_i[31]), .B(N0), .Z(N2) );
  GTECH_AND2 C21 ( .A(N354), .B(N275), .Z(N3) );
  GTECH_AND2 C22 ( .A(N414), .B(N202), .Z(N4) );
  GTECH_AND2 C24 ( .A(N321), .B(N136), .Z(N5) );
  GTECH_AND2 C28 ( .A(N2), .B(N3), .Z(N6) );
  GTECH_AND2 C29 ( .A(N4), .B(N206), .Z(N7) );
  GTECH_AND2 C30 ( .A(N5), .B(N138), .Z(N8) );
  GTECH_AND2 C32 ( .A(N6), .B(N7), .Z(N9) );
  GTECH_AND2 C33 ( .A(N8), .B(N141), .Z(N10) );
  GTECH_AND2 C34 ( .A(N9), .B(N10), .Z(N11) );
  GTECH_AND2 C35 ( .A(N11), .B(N1), .Z(N12) );
  GTECH_AND2 C52 ( .A(inp_i[30]), .B(N0), .Z(N13) );
  GTECH_AND2 C60 ( .A(N13), .B(N3), .Z(N14) );
  GTECH_AND2 C64 ( .A(N14), .B(N7), .Z(N15) );
  GTECH_AND2 C66 ( .A(N15), .B(N10), .Z(N16) );
  GTECH_AND2 C67 ( .A(N16), .B(N1), .Z(N17) );
  GTECH_AND2 C84 ( .A(inp_i[29]), .B(N0), .Z(N18) );
  GTECH_AND2 C92 ( .A(N18), .B(N3), .Z(N19) );
  GTECH_AND2 C96 ( .A(N19), .B(N7), .Z(N20) );
  GTECH_AND2 C98 ( .A(N20), .B(N10), .Z(N21) );
  GTECH_AND2 C99 ( .A(N21), .B(N1), .Z(N22) );
  GTECH_AND2 C116 ( .A(inp_i[28]), .B(N0), .Z(N23) );
  GTECH_AND2 C124 ( .A(N23), .B(N3), .Z(N24) );
  GTECH_AND2 C128 ( .A(N24), .B(N7), .Z(N25) );
  GTECH_AND2 C130 ( .A(N25), .B(N10), .Z(N26) );
  GTECH_AND2 C131 ( .A(N26), .B(N1), .Z(N27) );
  GTECH_AND2 C148 ( .A(inp_i[27]), .B(N0), .Z(N28) );
  GTECH_AND2 C156 ( .A(N28), .B(N3), .Z(N29) );
  GTECH_AND2 C160 ( .A(N29), .B(N7), .Z(N30) );
  GTECH_AND2 C162 ( .A(N30), .B(N10), .Z(N31) );
  GTECH_AND2 C163 ( .A(N31), .B(N1), .Z(N32) );
  GTECH_AND2 C180 ( .A(inp_i[26]), .B(N0), .Z(N33) );
  GTECH_AND2 C188 ( .A(N33), .B(N3), .Z(N34) );
  GTECH_AND2 C192 ( .A(N34), .B(N7), .Z(N35) );
  GTECH_AND2 C194 ( .A(N35), .B(N10), .Z(N36) );
  GTECH_AND2 C195 ( .A(N36), .B(N1), .Z(N37) );
  GTECH_AND2 C212 ( .A(inp_i[25]), .B(N0), .Z(N38) );
  GTECH_AND2 C220 ( .A(N38), .B(N3), .Z(N39) );
  GTECH_AND2 C224 ( .A(N39), .B(N7), .Z(N40) );
  GTECH_AND2 C226 ( .A(N40), .B(N10), .Z(N41) );
  GTECH_AND2 C227 ( .A(N41), .B(N1), .Z(N42) );
  GTECH_AND2 C244 ( .A(inp_i[24]), .B(N0), .Z(N43) );
  GTECH_AND2 C252 ( .A(N43), .B(N3), .Z(N44) );
  GTECH_AND2 C256 ( .A(N44), .B(N7), .Z(N45) );
  GTECH_AND2 C258 ( .A(N45), .B(N10), .Z(N46) );
  GTECH_AND2 C259 ( .A(N46), .B(N1), .Z(N47) );
  GTECH_AND2 C276 ( .A(inp_i[23]), .B(N0), .Z(N48) );
  GTECH_AND2 C284 ( .A(N48), .B(N3), .Z(N49) );
  GTECH_AND2 C288 ( .A(N49), .B(N7), .Z(N50) );
  GTECH_AND2 C290 ( .A(N50), .B(N10), .Z(N51) );
  GTECH_AND2 C291 ( .A(N51), .B(N1), .Z(N52) );
  GTECH_AND2 C308 ( .A(inp_i[22]), .B(N0), .Z(N53) );
  GTECH_AND2 C316 ( .A(N53), .B(N3), .Z(N54) );
  GTECH_AND2 C320 ( .A(N54), .B(N7), .Z(N55) );
  GTECH_AND2 C322 ( .A(N55), .B(N10), .Z(N56) );
  GTECH_AND2 C323 ( .A(N56), .B(N1), .Z(N57) );
  GTECH_AND2 C340 ( .A(inp_i[21]), .B(N0), .Z(N58) );
  GTECH_AND2 C348 ( .A(N58), .B(N3), .Z(N59) );
  GTECH_AND2 C352 ( .A(N59), .B(N7), .Z(N60) );
  GTECH_AND2 C354 ( .A(N60), .B(N10), .Z(N61) );
  GTECH_AND2 C355 ( .A(N61), .B(N1), .Z(N62) );
  GTECH_AND2 C372 ( .A(inp_i[20]), .B(N0), .Z(N63) );
  GTECH_AND2 C380 ( .A(N63), .B(N3), .Z(N64) );
  GTECH_AND2 C384 ( .A(N64), .B(N7), .Z(N65) );
  GTECH_AND2 C386 ( .A(N65), .B(N10), .Z(N66) );
  GTECH_AND2 C387 ( .A(N66), .B(N1), .Z(N67) );
  GTECH_AND2 C404 ( .A(inp_i[19]), .B(N0), .Z(N68) );
  GTECH_AND2 C412 ( .A(N68), .B(N3), .Z(N69) );
  GTECH_AND2 C416 ( .A(N69), .B(N7), .Z(N70) );
  GTECH_AND2 C418 ( .A(N70), .B(N10), .Z(N71) );
  GTECH_AND2 C419 ( .A(N71), .B(N1), .Z(N72) );
  GTECH_AND2 C436 ( .A(inp_i[18]), .B(N0), .Z(N73) );
  GTECH_AND2 C444 ( .A(N73), .B(N3), .Z(N74) );
  GTECH_AND2 C448 ( .A(N74), .B(N7), .Z(N75) );
  GTECH_AND2 C450 ( .A(N75), .B(N10), .Z(N76) );
  GTECH_AND2 C451 ( .A(N76), .B(N1), .Z(N77) );
  GTECH_AND2 C468 ( .A(inp_i[17]), .B(N0), .Z(N78) );
  GTECH_AND2 C476 ( .A(N78), .B(N3), .Z(N79) );
  GTECH_AND2 C480 ( .A(N79), .B(N7), .Z(N80) );
  GTECH_AND2 C482 ( .A(N80), .B(N10), .Z(N81) );
  GTECH_AND2 C483 ( .A(N81), .B(N1), .Z(N82) );
  GTECH_AND2 C500 ( .A(inp_i[16]), .B(N0), .Z(N83) );
  GTECH_AND2 C508 ( .A(N83), .B(N3), .Z(N84) );
  GTECH_AND2 C512 ( .A(N84), .B(N7), .Z(N85) );
  GTECH_AND2 C514 ( .A(N85), .B(N10), .Z(N86) );
  GTECH_AND2 C515 ( .A(N86), .B(N1), .Z(N87) );
  GTECH_AND2 C538 ( .A(inp_i[31]), .B(N89), .Z(N90) );
  GTECH_AND2 C539 ( .A(N353), .B(N273), .Z(N91) );
  GTECH_AND2 C540 ( .A(N274), .B(N198), .Z(N92) );
  GTECH_AND2 C542 ( .A(N201), .B(N136), .Z(N93) );
  GTECH_AND2 C546 ( .A(N90), .B(N91), .Z(N94) );
  GTECH_AND2 C547 ( .A(N92), .B(N204), .Z(N95) );
  GTECH_AND2 C548 ( .A(N93), .B(N138), .Z(N96) );
  GTECH_AND2 C550 ( .A(N94), .B(N95), .Z(N97) );
  GTECH_AND2 C551 ( .A(N96), .B(N141), .Z(N98) );
  GTECH_AND2 C552 ( .A(N97), .B(N98), .Z(N99) );
  GTECH_AND2 C553 ( .A(N99), .B(N1), .Z(N100) );
  GTECH_AND2 C570 ( .A(inp_i[30]), .B(N89), .Z(N101) );
  GTECH_AND2 C578 ( .A(N101), .B(N91), .Z(N102) );
  GTECH_AND2 C582 ( .A(N102), .B(N95), .Z(N103) );
  GTECH_AND2 C584 ( .A(N103), .B(N98), .Z(N104) );
  GTECH_AND2 C585 ( .A(N104), .B(N1), .Z(N105) );
  GTECH_AND2 C602 ( .A(inp_i[29]), .B(N89), .Z(N106) );
  GTECH_AND2 C610 ( .A(N106), .B(N91), .Z(N107) );
  GTECH_AND2 C614 ( .A(N107), .B(N95), .Z(N108) );
  GTECH_AND2 C616 ( .A(N108), .B(N98), .Z(N109) );
  GTECH_AND2 C617 ( .A(N109), .B(N1), .Z(N110) );
  GTECH_AND2 C634 ( .A(inp_i[28]), .B(N89), .Z(N111) );
  GTECH_AND2 C642 ( .A(N111), .B(N91), .Z(N112) );
  GTECH_AND2 C646 ( .A(N112), .B(N95), .Z(N113) );
  GTECH_AND2 C648 ( .A(N113), .B(N98), .Z(N114) );
  GTECH_AND2 C649 ( .A(N114), .B(N1), .Z(N115) );
  GTECH_AND2 C666 ( .A(inp_i[27]), .B(N89), .Z(N116) );
  GTECH_AND2 C674 ( .A(N116), .B(N91), .Z(N117) );
  GTECH_AND2 C678 ( .A(N117), .B(N95), .Z(N118) );
  GTECH_AND2 C680 ( .A(N118), .B(N98), .Z(N119) );
  GTECH_AND2 C681 ( .A(N119), .B(N1), .Z(N120) );
  GTECH_AND2 C698 ( .A(inp_i[26]), .B(N89), .Z(N121) );
  GTECH_AND2 C706 ( .A(N121), .B(N91), .Z(N122) );
  GTECH_AND2 C710 ( .A(N122), .B(N95), .Z(N123) );
  GTECH_AND2 C712 ( .A(N123), .B(N98), .Z(N124) );
  GTECH_AND2 C713 ( .A(N124), .B(N1), .Z(N125) );
  GTECH_AND2 C730 ( .A(inp_i[25]), .B(N89), .Z(N126) );
  GTECH_AND2 C738 ( .A(N126), .B(N91), .Z(N127) );
  GTECH_AND2 C742 ( .A(N127), .B(N95), .Z(N128) );
  GTECH_AND2 C744 ( .A(N128), .B(N98), .Z(N129) );
  GTECH_AND2 C745 ( .A(N129), .B(N1), .Z(N130) );
  GTECH_AND2 C762 ( .A(inp_i[24]), .B(N89), .Z(N131) );
  GTECH_AND2 C770 ( .A(N131), .B(N91), .Z(N132) );
  GTECH_AND2 C774 ( .A(N132), .B(N95), .Z(N133) );
  GTECH_AND2 C776 ( .A(N133), .B(N98), .Z(N134) );
  GTECH_AND2 C777 ( .A(N134), .B(N1), .Z(N135) );
  GTECH_AND2 C786 ( .A(inp_i[15]), .B(N136), .Z(N137) );
  GTECH_AND2 C787 ( .A(N391), .B(N322), .Z(N138) );
  GTECH_AND2 C788 ( .A(N430), .B(N242), .Z(N139) );
  GTECH_AND2 C790 ( .A(N137), .B(N138), .Z(N140) );
  GTECH_AND2 C791 ( .A(N139), .B(N244), .Z(N141) );
  GTECH_AND2 C792 ( .A(N140), .B(N141), .Z(N142) );
  GTECH_AND2 C793 ( .A(N142), .B(N1), .Z(N143) );
  GTECH_AND2 C802 ( .A(inp_i[14]), .B(N136), .Z(N144) );
  GTECH_AND2 C806 ( .A(N144), .B(N138), .Z(N145) );
  GTECH_AND2 C808 ( .A(N145), .B(N141), .Z(N146) );
  GTECH_AND2 C809 ( .A(N146), .B(N1), .Z(N147) );
  GTECH_AND2 C818 ( .A(inp_i[13]), .B(N136), .Z(N148) );
  GTECH_AND2 C822 ( .A(N148), .B(N138), .Z(N149) );
  GTECH_AND2 C824 ( .A(N149), .B(N141), .Z(N150) );
  GTECH_AND2 C825 ( .A(N150), .B(N1), .Z(N151) );
  GTECH_AND2 C834 ( .A(inp_i[12]), .B(N136), .Z(N152) );
  GTECH_AND2 C838 ( .A(N152), .B(N138), .Z(N153) );
  GTECH_AND2 C840 ( .A(N153), .B(N141), .Z(N154) );
  GTECH_AND2 C841 ( .A(N154), .B(N1), .Z(N155) );
  GTECH_AND2 C850 ( .A(inp_i[11]), .B(N136), .Z(N156) );
  GTECH_AND2 C854 ( .A(N156), .B(N138), .Z(N157) );
  GTECH_AND2 C856 ( .A(N157), .B(N141), .Z(N158) );
  GTECH_AND2 C857 ( .A(N158), .B(N1), .Z(N159) );
  GTECH_AND2 C866 ( .A(inp_i[10]), .B(N136), .Z(N160) );
  GTECH_AND2 C870 ( .A(N160), .B(N138), .Z(N161) );
  GTECH_AND2 C872 ( .A(N161), .B(N141), .Z(N162) );
  GTECH_AND2 C873 ( .A(N162), .B(N1), .Z(N163) );
  GTECH_AND2 C882 ( .A(inp_i[9]), .B(N136), .Z(N164) );
  GTECH_AND2 C886 ( .A(N164), .B(N138), .Z(N165) );
  GTECH_AND2 C888 ( .A(N165), .B(N141), .Z(N166) );
  GTECH_AND2 C889 ( .A(N166), .B(N1), .Z(N167) );
  GTECH_AND2 C898 ( .A(inp_i[8]), .B(N136), .Z(N168) );
  GTECH_AND2 C902 ( .A(N168), .B(N138), .Z(N169) );
  GTECH_AND2 C904 ( .A(N169), .B(N141), .Z(N170) );
  GTECH_AND2 C905 ( .A(N170), .B(N1), .Z(N171) );
  GTECH_AND2 C928 ( .A(inp_i[31]), .B(N173), .Z(N174) );
  GTECH_AND2 C929 ( .A(N352), .B(N271), .Z(N175) );
  GTECH_AND2 C930 ( .A(N272), .B(N198), .Z(N176) );
  GTECH_AND2 C936 ( .A(N174), .B(N175), .Z(N177) );
  GTECH_AND2 C937 ( .A(N176), .B(N204), .Z(N178) );
  GTECH_AND2 C940 ( .A(N177), .B(N178), .Z(N179) );
  GTECH_AND2 C941 ( .A(N209), .B(N210), .Z(N180) );
  GTECH_AND2 C942 ( .A(N179), .B(N180), .Z(N181) );
  GTECH_AND2 C943 ( .A(N181), .B(N1), .Z(N182) );
  GTECH_AND2 C960 ( .A(inp_i[30]), .B(N173), .Z(N183) );
  GTECH_AND2 C968 ( .A(N183), .B(N175), .Z(N184) );
  GTECH_AND2 C972 ( .A(N184), .B(N178), .Z(N185) );
  GTECH_AND2 C974 ( .A(N185), .B(N180), .Z(N186) );
  GTECH_AND2 C975 ( .A(N186), .B(N1), .Z(N187) );
  GTECH_AND2 C992 ( .A(inp_i[29]), .B(N173), .Z(N188) );
  GTECH_AND2 C1000 ( .A(N188), .B(N175), .Z(N189) );
  GTECH_AND2 C1004 ( .A(N189), .B(N178), .Z(N190) );
  GTECH_AND2 C1006 ( .A(N190), .B(N180), .Z(N191) );
  GTECH_AND2 C1007 ( .A(N191), .B(N1), .Z(N192) );
  GTECH_AND2 C1024 ( .A(inp_i[28]), .B(N173), .Z(N193) );
  GTECH_AND2 C1032 ( .A(N193), .B(N175), .Z(N194) );
  GTECH_AND2 C1036 ( .A(N194), .B(N178), .Z(N195) );
  GTECH_AND2 C1038 ( .A(N195), .B(N180), .Z(N196) );
  GTECH_AND2 C1039 ( .A(N196), .B(N1), .Z(N197) );
  GTECH_AND2 C1052 ( .A(inp_i[23]), .B(N198), .Z(N203) );
  GTECH_AND2 C1053 ( .A(N199), .B(N200), .Z(N204) );
  GTECH_AND2 C1054 ( .A(N201), .B(N202), .Z(N205) );
  GTECH_AND2 C1055 ( .A(N415), .B(N320), .Z(N206) );
  GTECH_AND2 C1056 ( .A(N321), .B(N242), .Z(N207) );
  GTECH_AND2 C1058 ( .A(N203), .B(N204), .Z(N208) );
  GTECH_AND2 C1059 ( .A(N205), .B(N206), .Z(N209) );
  GTECH_AND2 C1060 ( .A(N207), .B(N244), .Z(N210) );
  GTECH_AND2 C1061 ( .A(N208), .B(N209), .Z(N211) );
  GTECH_AND2 C1062 ( .A(N210), .B(N1), .Z(N212) );
  GTECH_AND2 C1063 ( .A(N211), .B(N212), .Z(N213) );
  GTECH_AND2 C1076 ( .A(inp_i[22]), .B(N198), .Z(N214) );
  GTECH_AND2 C1082 ( .A(N214), .B(N204), .Z(N215) );
  GTECH_AND2 C1085 ( .A(N215), .B(N209), .Z(N216) );
  GTECH_AND2 C1087 ( .A(N216), .B(N212), .Z(N217) );
  GTECH_AND2 C1100 ( .A(inp_i[21]), .B(N198), .Z(N218) );
  GTECH_AND2 C1106 ( .A(N218), .B(N204), .Z(N219) );
  GTECH_AND2 C1109 ( .A(N219), .B(N209), .Z(N220) );
  GTECH_AND2 C1111 ( .A(N220), .B(N212), .Z(N221) );
  GTECH_AND2 C1124 ( .A(inp_i[20]), .B(N198), .Z(N222) );
  GTECH_AND2 C1130 ( .A(N222), .B(N204), .Z(N223) );
  GTECH_AND2 C1133 ( .A(N223), .B(N209), .Z(N224) );
  GTECH_AND2 C1135 ( .A(N224), .B(N212), .Z(N225) );
  GTECH_AND2 C1144 ( .A(inp_i[15]), .B(N202), .Z(N226) );
  GTECH_AND2 C1148 ( .A(N226), .B(N206), .Z(N227) );
  GTECH_AND2 C1150 ( .A(N227), .B(N210), .Z(N228) );
  GTECH_AND2 C1151 ( .A(N228), .B(N1), .Z(N229) );
  GTECH_AND2 C1160 ( .A(inp_i[14]), .B(N202), .Z(N230) );
  GTECH_AND2 C1164 ( .A(N230), .B(N206), .Z(N231) );
  GTECH_AND2 C1166 ( .A(N231), .B(N210), .Z(N232) );
  GTECH_AND2 C1167 ( .A(N232), .B(N1), .Z(N233) );
  GTECH_AND2 C1176 ( .A(inp_i[13]), .B(N202), .Z(N234) );
  GTECH_AND2 C1180 ( .A(N234), .B(N206), .Z(N235) );
  GTECH_AND2 C1182 ( .A(N235), .B(N210), .Z(N236) );
  GTECH_AND2 C1183 ( .A(N236), .B(N1), .Z(N237) );
  GTECH_AND2 C1192 ( .A(inp_i[12]), .B(N202), .Z(N238) );
  GTECH_AND2 C1196 ( .A(N238), .B(N206), .Z(N239) );
  GTECH_AND2 C1198 ( .A(N239), .B(N210), .Z(N240) );
  GTECH_AND2 C1199 ( .A(N240), .B(N1), .Z(N241) );
  GTECH_AND2 C1204 ( .A(inp_i[7]), .B(N242), .Z(N243) );
  GTECH_AND2 C1205 ( .A(N404), .B(N336), .Z(N244) );
  GTECH_AND2 C1206 ( .A(N243), .B(N244), .Z(N245) );
  GTECH_AND2 C1207 ( .A(N245), .B(N1), .Z(N246) );
  GTECH_AND2 C1212 ( .A(inp_i[6]), .B(N242), .Z(N247) );
  GTECH_AND2 C1214 ( .A(N247), .B(N244), .Z(N248) );
  GTECH_AND2 C1215 ( .A(N248), .B(N1), .Z(N249) );
  GTECH_AND2 C1220 ( .A(inp_i[5]), .B(N242), .Z(N250) );
  GTECH_AND2 C1222 ( .A(N250), .B(N244), .Z(N251) );
  GTECH_AND2 C1223 ( .A(N251), .B(N1), .Z(N252) );
  GTECH_AND2 C1228 ( .A(inp_i[4]), .B(N242), .Z(N253) );
  GTECH_AND2 C1230 ( .A(N253), .B(N244), .Z(N254) );
  GTECH_AND2 C1231 ( .A(N254), .B(N1), .Z(N255) );
  GTECH_AND2 C1254 ( .A(inp_i[31]), .B(N257), .Z(N258) );
  GTECH_AND2 C1255 ( .A(N351), .B(N271), .Z(N259) );
  GTECH_AND2 C1262 ( .A(N258), .B(N259), .Z(N260) );
  GTECH_AND2 C1263 ( .A(N277), .B(N278), .Z(N261) );
  GTECH_AND2 C1266 ( .A(N260), .B(N261), .Z(N262) );
  GTECH_AND2 C1267 ( .A(N293), .B(N294), .Z(N263) );
  GTECH_AND2 C1268 ( .A(N262), .B(N263), .Z(N264) );
  GTECH_AND2 C1269 ( .A(N264), .B(N1), .Z(N265) );
  GTECH_AND2 C1286 ( .A(inp_i[30]), .B(N257), .Z(N266) );
  GTECH_AND2 C1294 ( .A(N266), .B(N259), .Z(N267) );
  GTECH_AND2 C1298 ( .A(N267), .B(N261), .Z(N268) );
  GTECH_AND2 C1300 ( .A(N268), .B(N263), .Z(N269) );
  GTECH_AND2 C1301 ( .A(N269), .B(N1), .Z(N270) );
  GTECH_AND2 C1316 ( .A(inp_i[27]), .B(N271), .Z(N276) );
  GTECH_AND2 C1317 ( .A(N272), .B(N273), .Z(N277) );
  GTECH_AND2 C1318 ( .A(N274), .B(N200), .Z(N278) );
  GTECH_AND2 C1319 ( .A(N201), .B(N275), .Z(N279) );
  GTECH_AND2 C1320 ( .A(N414), .B(N320), .Z(N280) );
  GTECH_AND2 C1323 ( .A(N276), .B(N277), .Z(N281) );
  GTECH_AND2 C1324 ( .A(N278), .B(N279), .Z(N282) );
  GTECH_AND2 C1325 ( .A(N280), .B(N324), .Z(N283) );
  GTECH_AND2 C1327 ( .A(N281), .B(N282), .Z(N284) );
  GTECH_AND2 C1328 ( .A(N283), .B(N305), .Z(N285) );
  GTECH_AND2 C1329 ( .A(N284), .B(N285), .Z(N286) );
  GTECH_AND2 C1344 ( .A(inp_i[26]), .B(N271), .Z(N287) );
  GTECH_AND2 C1351 ( .A(N287), .B(N277), .Z(N288) );
  GTECH_AND2 C1355 ( .A(N288), .B(N282), .Z(N289) );
  GTECH_AND2 C1357 ( .A(N289), .B(N285), .Z(N290) );
  GTECH_AND2 C1370 ( .A(inp_i[23]), .B(N273), .Z(N291) );
  GTECH_AND2 C1376 ( .A(N291), .B(N278), .Z(N292) );
  GTECH_AND2 C1377 ( .A(N279), .B(N280), .Z(N293) );
  GTECH_AND2 C1378 ( .A(N324), .B(N303), .Z(N294) );
  GTECH_AND2 C1379 ( .A(N292), .B(N293), .Z(N295) );
  GTECH_AND2 C1380 ( .A(N294), .B(N1), .Z(N296) );
  GTECH_AND2 C1381 ( .A(N295), .B(N296), .Z(N297) );
  GTECH_AND2 C1394 ( .A(inp_i[22]), .B(N273), .Z(N298) );
  GTECH_AND2 C1400 ( .A(N298), .B(N278), .Z(N299) );
  GTECH_AND2 C1403 ( .A(N299), .B(N293), .Z(N300) );
  GTECH_AND2 C1405 ( .A(N300), .B(N296), .Z(N301) );
  GTECH_AND2 C1416 ( .A(inp_i[19]), .B(N200), .Z(N302) );
  GTECH_AND2 C1420 ( .A(N430), .B(N336), .Z(N303) );
  GTECH_AND2 C1421 ( .A(N302), .B(N279), .Z(N304) );
  GTECH_AND2 C1423 ( .A(N303), .B(N1), .Z(N305) );
  GTECH_AND2 C1424 ( .A(N304), .B(N283), .Z(N306) );
  GTECH_AND2 C1425 ( .A(N306), .B(N305), .Z(N307) );
  GTECH_AND2 C1436 ( .A(inp_i[18]), .B(N200), .Z(N308) );
  GTECH_AND2 C1441 ( .A(N308), .B(N279), .Z(N309) );
  GTECH_AND2 C1444 ( .A(N309), .B(N283), .Z(N310) );
  GTECH_AND2 C1445 ( .A(N310), .B(N305), .Z(N311) );
  GTECH_AND2 C1454 ( .A(inp_i[15]), .B(N275), .Z(N312) );
  GTECH_AND2 C1458 ( .A(N312), .B(N280), .Z(N313) );
  GTECH_AND2 C1460 ( .A(N313), .B(N294), .Z(N314) );
  GTECH_AND2 C1461 ( .A(N314), .B(N1), .Z(N315) );
  GTECH_AND2 C1470 ( .A(inp_i[14]), .B(N275), .Z(N316) );
  GTECH_AND2 C1474 ( .A(N316), .B(N280), .Z(N317) );
  GTECH_AND2 C1476 ( .A(N317), .B(N294), .Z(N318) );
  GTECH_AND2 C1477 ( .A(N318), .B(N1), .Z(N319) );
  GTECH_AND2 C1484 ( .A(inp_i[11]), .B(N320), .Z(N323) );
  GTECH_AND2 C1485 ( .A(N321), .B(N322), .Z(N324) );
  GTECH_AND2 C1487 ( .A(N323), .B(N324), .Z(N325) );
  GTECH_AND2 C1489 ( .A(N325), .B(N305), .Z(N326) );
  GTECH_AND2 C1496 ( .A(inp_i[10]), .B(N320), .Z(N327) );
  GTECH_AND2 C1499 ( .A(N327), .B(N324), .Z(N328) );
  GTECH_AND2 C1501 ( .A(N328), .B(N305), .Z(N329) );
  GTECH_AND2 C1506 ( .A(inp_i[7]), .B(N322), .Z(N330) );
  GTECH_AND2 C1508 ( .A(N330), .B(N303), .Z(N331) );
  GTECH_AND2 C1509 ( .A(N331), .B(N1), .Z(N332) );
  GTECH_AND2 C1514 ( .A(inp_i[6]), .B(N322), .Z(N333) );
  GTECH_AND2 C1516 ( .A(N333), .B(N303), .Z(N334) );
  GTECH_AND2 C1517 ( .A(N334), .B(N1), .Z(N335) );
  GTECH_AND2 C1520 ( .A(inp_i[3]), .B(N336), .Z(N337) );
  GTECH_AND2 C1521 ( .A(N337), .B(N1), .Z(N338) );
  GTECH_AND2 C1524 ( .A(inp_i[2]), .B(N336), .Z(N339) );
  GTECH_AND2 C1525 ( .A(N339), .B(N1), .Z(N340) );
  GTECH_AND2 C1548 ( .A(inp_i[31]), .B(N342), .Z(N343) );
  GTECH_AND2 C1549 ( .A(N351), .B(N352), .Z(N344) );
  GTECH_AND2 C1556 ( .A(N343), .B(N344), .Z(N345) );
  GTECH_AND2 C1557 ( .A(N367), .B(N368), .Z(N346) );
  GTECH_AND2 C1560 ( .A(N345), .B(N346), .Z(N347) );
  GTECH_AND2 C1561 ( .A(N386), .B(N387), .Z(N348) );
  GTECH_AND2 C1562 ( .A(N347), .B(N348), .Z(N349) );
  GTECH_AND2 C1563 ( .A(N349), .B(N1), .Z(N350) );
  GTECH_AND2 C1579 ( .A(inp_i[29]), .B(N351), .Z(N355) );
  GTECH_AND2 C1580 ( .A(N352), .B(N272), .Z(N356) );
  GTECH_AND2 C1581 ( .A(N353), .B(N274), .Z(N357) );
  GTECH_AND2 C1582 ( .A(N199), .B(N201), .Z(N358) );
  GTECH_AND2 C1583 ( .A(N354), .B(N414), .Z(N359) );
  GTECH_AND2 C1587 ( .A(N355), .B(N356), .Z(N360) );
  GTECH_AND2 C1588 ( .A(N357), .B(N358), .Z(N361) );
  GTECH_AND2 C1589 ( .A(N359), .B(N417), .Z(N362) );
  GTECH_AND2 C1591 ( .A(N360), .B(N361), .Z(N363) );
  GTECH_AND2 C1592 ( .A(N362), .B(N395), .Z(N364) );
  GTECH_AND2 C1593 ( .A(N363), .B(N364), .Z(N365) );
  GTECH_AND2 C1608 ( .A(inp_i[27]), .B(N352), .Z(N366) );
  GTECH_AND2 C1609 ( .A(N272), .B(N353), .Z(N367) );
  GTECH_AND2 C1610 ( .A(N274), .B(N199), .Z(N368) );
  GTECH_AND2 C1611 ( .A(N201), .B(N354), .Z(N369) );
  GTECH_AND2 C1612 ( .A(N414), .B(N415), .Z(N370) );
  GTECH_AND2 C1615 ( .A(N366), .B(N367), .Z(N371) );
  GTECH_AND2 C1616 ( .A(N368), .B(N369), .Z(N372) );
  GTECH_AND2 C1617 ( .A(N370), .B(N421), .Z(N373) );
  GTECH_AND2 C1619 ( .A(N371), .B(N372), .Z(N374) );
  GTECH_AND2 C1620 ( .A(N373), .B(N401), .Z(N375) );
  GTECH_AND2 C1621 ( .A(N374), .B(N375), .Z(N376) );
  GTECH_AND2 C1635 ( .A(inp_i[25]), .B(N272), .Z(N377) );
  GTECH_AND2 C1642 ( .A(N377), .B(N357), .Z(N378) );
  GTECH_AND2 C1643 ( .A(N358), .B(N359), .Z(N379) );
  GTECH_AND2 C1644 ( .A(N417), .B(N393), .Z(N380) );
  GTECH_AND2 C1645 ( .A(N378), .B(N379), .Z(N381) );
  GTECH_AND2 C1646 ( .A(N380), .B(N406), .Z(N382) );
  GTECH_AND2 C1647 ( .A(N381), .B(N382), .Z(N383) );
  GTECH_AND2 C1660 ( .A(inp_i[23]), .B(N353), .Z(N384) );
  GTECH_AND2 C1666 ( .A(N384), .B(N368), .Z(N385) );
  GTECH_AND2 C1667 ( .A(N369), .B(N370), .Z(N386) );
  GTECH_AND2 C1668 ( .A(N421), .B(N399), .Z(N387) );
  GTECH_AND2 C1669 ( .A(N385), .B(N386), .Z(N388) );
  GTECH_AND2 C1670 ( .A(N387), .B(N1), .Z(N389) );
  GTECH_AND2 C1671 ( .A(N388), .B(N389), .Z(N390) );
  GTECH_AND2 C1683 ( .A(inp_i[21]), .B(N274), .Z(N392) );
  GTECH_AND2 C1687 ( .A(N391), .B(N430), .Z(N393) );
  GTECH_AND2 C1689 ( .A(N392), .B(N358), .Z(N394) );
  GTECH_AND2 C1691 ( .A(N393), .B(N406), .Z(N395) );
  GTECH_AND2 C1692 ( .A(N394), .B(N362), .Z(N396) );
  GTECH_AND2 C1693 ( .A(N396), .B(N395), .Z(N397) );
  GTECH_AND2 C1704 ( .A(inp_i[19]), .B(N199), .Z(N398) );
  GTECH_AND2 C1708 ( .A(N430), .B(N404), .Z(N399) );
  GTECH_AND2 C1709 ( .A(N398), .B(N369), .Z(N400) );
  GTECH_AND2 C1711 ( .A(N399), .B(N1), .Z(N401) );
  GTECH_AND2 C1712 ( .A(N400), .B(N373), .Z(N402) );
  GTECH_AND2 C1713 ( .A(N402), .B(N401), .Z(N403) );
  GTECH_AND2 C1723 ( .A(inp_i[17]), .B(N201), .Z(N405) );
  GTECH_AND2 C1727 ( .A(N404), .B(N1), .Z(N406) );
  GTECH_AND2 C1728 ( .A(N405), .B(N359), .Z(N407) );
  GTECH_AND2 C1730 ( .A(N407), .B(N380), .Z(N408) );
  GTECH_AND2 C1731 ( .A(N408), .B(N406), .Z(N409) );
  GTECH_AND2 C1740 ( .A(inp_i[15]), .B(N354), .Z(N410) );
  GTECH_AND2 C1744 ( .A(N410), .B(N370), .Z(N411) );
  GTECH_AND2 C1746 ( .A(N411), .B(N387), .Z(N412) );
  GTECH_AND2 C1747 ( .A(N412), .B(N1), .Z(N413) );
  GTECH_AND2 C1755 ( .A(inp_i[13]), .B(N414), .Z(N416) );
  GTECH_AND2 C1756 ( .A(N415), .B(N321), .Z(N417) );
  GTECH_AND2 C1759 ( .A(N416), .B(N417), .Z(N418) );
  GTECH_AND2 C1761 ( .A(N418), .B(N395), .Z(N419) );
  GTECH_AND2 C1768 ( .A(inp_i[11]), .B(N415), .Z(N420) );
  GTECH_AND2 C1769 ( .A(N321), .B(N391), .Z(N421) );
  GTECH_AND2 C1771 ( .A(N420), .B(N421), .Z(N422) );
  GTECH_AND2 C1773 ( .A(N422), .B(N401), .Z(N423) );
  GTECH_AND2 C1779 ( .A(inp_i[9]), .B(N321), .Z(N424) );
  GTECH_AND2 C1782 ( .A(N424), .B(N393), .Z(N425) );
  GTECH_AND2 C1783 ( .A(N425), .B(N406), .Z(N426) );
  GTECH_AND2 C1788 ( .A(inp_i[7]), .B(N391), .Z(N427) );
  GTECH_AND2 C1790 ( .A(N427), .B(N399), .Z(N428) );
  GTECH_AND2 C1791 ( .A(N428), .B(N1), .Z(N429) );
  GTECH_AND2 C1795 ( .A(inp_i[5]), .B(N430), .Z(N431) );
  GTECH_AND2 C1797 ( .A(N431), .B(N406), .Z(N432) );
  GTECH_AND2 C1800 ( .A(inp_i[3]), .B(N404), .Z(N433) );
  GTECH_AND2 C1801 ( .A(N433), .B(N1), .Z(N434) );
  GTECH_AND2 C1803 ( .A(inp_i[1]), .B(N1), .Z(N435) );
  GTECH_OR2 C1816 ( .A(inp_i[30]), .B(inp_i[31]), .Z(N437) );
  GTECH_OR2 C1817 ( .A(inp_i[29]), .B(N437), .Z(N438) );
  GTECH_OR2 C1818 ( .A(inp_i[28]), .B(N438), .Z(N439) );
  GTECH_OR2 C1819 ( .A(inp_i[27]), .B(N439), .Z(N440) );
  GTECH_OR2 C1820 ( .A(inp_i[26]), .B(N440), .Z(N441) );
  GTECH_OR2 C1821 ( .A(inp_i[25]), .B(N441), .Z(N442) );
  GTECH_OR2 C1822 ( .A(inp_i[24]), .B(N442), .Z(N443) );
  GTECH_OR2 C1823 ( .A(inp_i[23]), .B(N443), .Z(N444) );
  GTECH_OR2 C1824 ( .A(inp_i[22]), .B(N444), .Z(N445) );
  GTECH_OR2 C1825 ( .A(inp_i[21]), .B(N445), .Z(N446) );
  GTECH_OR2 C1826 ( .A(inp_i[20]), .B(N446), .Z(N447) );
  GTECH_OR2 C1827 ( .A(inp_i[19]), .B(N447), .Z(N448) );
  GTECH_OR2 C1828 ( .A(inp_i[18]), .B(N448), .Z(N449) );
  GTECH_OR2 C1829 ( .A(inp_i[17]), .B(N449), .Z(N450) );
  GTECH_OR2 C1830 ( .A(inp_i[16]), .B(N450), .Z(N451) );
  GTECH_OR2 C1831 ( .A(inp_i[15]), .B(N451), .Z(N452) );
  GTECH_OR2 C1832 ( .A(inp_i[14]), .B(N452), .Z(N453) );
  GTECH_OR2 C1833 ( .A(inp_i[13]), .B(N453), .Z(N454) );
  GTECH_OR2 C1834 ( .A(inp_i[12]), .B(N454), .Z(N455) );
  GTECH_OR2 C1835 ( .A(inp_i[11]), .B(N455), .Z(N456) );
  GTECH_OR2 C1836 ( .A(inp_i[10]), .B(N456), .Z(N457) );
  GTECH_OR2 C1837 ( .A(inp_i[9]), .B(N457), .Z(N458) );
  GTECH_OR2 C1838 ( .A(inp_i[8]), .B(N458), .Z(N459) );
  GTECH_OR2 C1839 ( .A(inp_i[7]), .B(N459), .Z(N460) );
  GTECH_OR2 C1840 ( .A(inp_i[6]), .B(N460), .Z(N461) );
  GTECH_OR2 C1841 ( .A(inp_i[5]), .B(N461), .Z(N462) );
  GTECH_OR2 C1842 ( .A(inp_i[4]), .B(N462), .Z(N463) );
  GTECH_OR2 C1843 ( .A(inp_i[3]), .B(N463), .Z(N464) );
  GTECH_OR2 C1844 ( .A(inp_i[2]), .B(N464), .Z(N465) );
  GTECH_OR2 C1845 ( .A(inp_i[1]), .B(N465), .Z(N466) );
  GTECH_OR2 C1846 ( .A(inp_i[0]), .B(N466), .Z(N467) );
  GTECH_NOT I_0 ( .A(N467), .Z(N468) );
  GTECH_NOT I_1 ( .A(N468), .Z(valid_o) );
  GTECH_NOT I_2 ( .A(inp_i[15]), .Z(N0) );
  GTECH_NOT I_3 ( .A(inp_i[0]), .Z(N1) );
  GTECH_OR2 C1852 ( .A(N12), .B(N482), .Z(N88) );
  GTECH_OR2 C1853 ( .A(N17), .B(N481), .Z(N482) );
  GTECH_OR2 C1854 ( .A(N22), .B(N480), .Z(N481) );
  GTECH_OR2 C1855 ( .A(N27), .B(N479), .Z(N480) );
  GTECH_OR2 C1856 ( .A(N32), .B(N478), .Z(N479) );
  GTECH_OR2 C1857 ( .A(N37), .B(N477), .Z(N478) );
  GTECH_OR2 C1858 ( .A(N42), .B(N476), .Z(N477) );
  GTECH_OR2 C1859 ( .A(N47), .B(N475), .Z(N476) );
  GTECH_OR2 C1860 ( .A(N52), .B(N474), .Z(N475) );
  GTECH_OR2 C1861 ( .A(N57), .B(N473), .Z(N474) );
  GTECH_OR2 C1862 ( .A(N62), .B(N472), .Z(N473) );
  GTECH_OR2 C1863 ( .A(N67), .B(N471), .Z(N472) );
  GTECH_OR2 C1864 ( .A(N72), .B(N470), .Z(N471) );
  GTECH_OR2 C1865 ( .A(N77), .B(N469), .Z(N470) );
  GTECH_OR2 C1866 ( .A(N82), .B(N87), .Z(N469) );
  GTECH_BUF B_0 ( .A(N88), .Z(out_o[4]) );
  GTECH_NOT I_4 ( .A(inp_i[23]), .Z(N89) );
  GTECH_NOT I_5 ( .A(inp_i[7]), .Z(N136) );
  GTECH_OR2 C1870 ( .A(N100), .B(N496), .Z(N172) );
  GTECH_OR2 C1871 ( .A(N105), .B(N495), .Z(N496) );
  GTECH_OR2 C1872 ( .A(N110), .B(N494), .Z(N495) );
  GTECH_OR2 C1873 ( .A(N115), .B(N493), .Z(N494) );
  GTECH_OR2 C1874 ( .A(N120), .B(N492), .Z(N493) );
  GTECH_OR2 C1875 ( .A(N125), .B(N491), .Z(N492) );
  GTECH_OR2 C1876 ( .A(N130), .B(N490), .Z(N491) );
  GTECH_OR2 C1877 ( .A(N135), .B(N489), .Z(N490) );
  GTECH_OR2 C1878 ( .A(N143), .B(N488), .Z(N489) );
  GTECH_OR2 C1879 ( .A(N147), .B(N487), .Z(N488) );
  GTECH_OR2 C1880 ( .A(N151), .B(N486), .Z(N487) );
  GTECH_OR2 C1881 ( .A(N155), .B(N485), .Z(N486) );
  GTECH_OR2 C1882 ( .A(N159), .B(N484), .Z(N485) );
  GTECH_OR2 C1883 ( .A(N163), .B(N483), .Z(N484) );
  GTECH_OR2 C1884 ( .A(N167), .B(N171), .Z(N483) );
  GTECH_BUF B_1 ( .A(N172), .Z(out_o[3]) );
  GTECH_NOT I_6 ( .A(inp_i[27]), .Z(N173) );
  GTECH_NOT I_7 ( .A(inp_i[19]), .Z(N198) );
  GTECH_NOT I_8 ( .A(inp_i[18]), .Z(N199) );
  GTECH_NOT I_9 ( .A(inp_i[17]), .Z(N200) );
  GTECH_NOT I_10 ( .A(inp_i[16]), .Z(N201) );
  GTECH_NOT I_11 ( .A(inp_i[11]), .Z(N202) );
  GTECH_NOT I_12 ( .A(inp_i[3]), .Z(N242) );
  GTECH_OR2 C1893 ( .A(N182), .B(N510), .Z(N256) );
  GTECH_OR2 C1894 ( .A(N187), .B(N509), .Z(N510) );
  GTECH_OR2 C1895 ( .A(N192), .B(N508), .Z(N509) );
  GTECH_OR2 C1896 ( .A(N197), .B(N507), .Z(N508) );
  GTECH_OR2 C1897 ( .A(N213), .B(N506), .Z(N507) );
  GTECH_OR2 C1898 ( .A(N217), .B(N505), .Z(N506) );
  GTECH_OR2 C1899 ( .A(N221), .B(N504), .Z(N505) );
  GTECH_OR2 C1900 ( .A(N225), .B(N503), .Z(N504) );
  GTECH_OR2 C1901 ( .A(N229), .B(N502), .Z(N503) );
  GTECH_OR2 C1902 ( .A(N233), .B(N501), .Z(N502) );
  GTECH_OR2 C1903 ( .A(N237), .B(N500), .Z(N501) );
  GTECH_OR2 C1904 ( .A(N241), .B(N499), .Z(N500) );
  GTECH_OR2 C1905 ( .A(N246), .B(N498), .Z(N499) );
  GTECH_OR2 C1906 ( .A(N249), .B(N497), .Z(N498) );
  GTECH_OR2 C1907 ( .A(N252), .B(N255), .Z(N497) );
  GTECH_BUF B_2 ( .A(N256), .Z(out_o[2]) );
  GTECH_NOT I_13 ( .A(inp_i[29]), .Z(N257) );
  GTECH_NOT I_14 ( .A(inp_i[25]), .Z(N271) );
  GTECH_NOT I_15 ( .A(inp_i[24]), .Z(N272) );
  GTECH_NOT I_16 ( .A(inp_i[21]), .Z(N273) );
  GTECH_NOT I_17 ( .A(inp_i[20]), .Z(N274) );
  GTECH_NOT I_18 ( .A(inp_i[13]), .Z(N275) );
  GTECH_NOT I_19 ( .A(inp_i[9]), .Z(N320) );
  GTECH_NOT I_20 ( .A(inp_i[8]), .Z(N321) );
  GTECH_NOT I_21 ( .A(inp_i[5]), .Z(N322) );
  GTECH_NOT I_22 ( .A(inp_i[1]), .Z(N336) );
  GTECH_OR2 C1919 ( .A(N265), .B(N524), .Z(N341) );
  GTECH_OR2 C1920 ( .A(N270), .B(N523), .Z(N524) );
  GTECH_OR2 C1921 ( .A(N286), .B(N522), .Z(N523) );
  GTECH_OR2 C1922 ( .A(N290), .B(N521), .Z(N522) );
  GTECH_OR2 C1923 ( .A(N297), .B(N520), .Z(N521) );
  GTECH_OR2 C1924 ( .A(N301), .B(N519), .Z(N520) );
  GTECH_OR2 C1925 ( .A(N307), .B(N518), .Z(N519) );
  GTECH_OR2 C1926 ( .A(N311), .B(N517), .Z(N518) );
  GTECH_OR2 C1927 ( .A(N315), .B(N516), .Z(N517) );
  GTECH_OR2 C1928 ( .A(N319), .B(N515), .Z(N516) );
  GTECH_OR2 C1929 ( .A(N326), .B(N514), .Z(N515) );
  GTECH_OR2 C1930 ( .A(N329), .B(N513), .Z(N514) );
  GTECH_OR2 C1931 ( .A(N332), .B(N512), .Z(N513) );
  GTECH_OR2 C1932 ( .A(N335), .B(N511), .Z(N512) );
  GTECH_OR2 C1933 ( .A(N338), .B(N340), .Z(N511) );
  GTECH_BUF B_3 ( .A(N341), .Z(out_o[1]) );
  GTECH_NOT I_23 ( .A(inp_i[30]), .Z(N342) );
  GTECH_NOT I_24 ( .A(inp_i[28]), .Z(N351) );
  GTECH_NOT I_25 ( .A(inp_i[26]), .Z(N352) );
  GTECH_NOT I_26 ( .A(inp_i[22]), .Z(N353) );
  GTECH_NOT I_27 ( .A(inp_i[14]), .Z(N354) );
  GTECH_NOT I_28 ( .A(inp_i[6]), .Z(N391) );
  GTECH_NOT I_29 ( .A(inp_i[2]), .Z(N404) );
  GTECH_NOT I_30 ( .A(inp_i[12]), .Z(N414) );
  GTECH_NOT I_31 ( .A(inp_i[10]), .Z(N415) );
  GTECH_NOT I_32 ( .A(inp_i[4]), .Z(N430) );
  GTECH_OR2 C1945 ( .A(N350), .B(N538), .Z(N436) );
  GTECH_OR2 C1946 ( .A(N365), .B(N537), .Z(N538) );
  GTECH_OR2 C1947 ( .A(N376), .B(N536), .Z(N537) );
  GTECH_OR2 C1948 ( .A(N383), .B(N535), .Z(N536) );
  GTECH_OR2 C1949 ( .A(N390), .B(N534), .Z(N535) );
  GTECH_OR2 C1950 ( .A(N397), .B(N533), .Z(N534) );
  GTECH_OR2 C1951 ( .A(N403), .B(N532), .Z(N533) );
  GTECH_OR2 C1952 ( .A(N409), .B(N531), .Z(N532) );
  GTECH_OR2 C1953 ( .A(N413), .B(N530), .Z(N531) );
  GTECH_OR2 C1954 ( .A(N419), .B(N529), .Z(N530) );
  GTECH_OR2 C1955 ( .A(N423), .B(N528), .Z(N529) );
  GTECH_OR2 C1956 ( .A(N426), .B(N527), .Z(N528) );
  GTECH_OR2 C1957 ( .A(N429), .B(N526), .Z(N527) );
  GTECH_OR2 C1958 ( .A(N432), .B(N525), .Z(N526) );
  GTECH_OR2 C1959 ( .A(N434), .B(N435), .Z(N525) );
  GTECH_BUF B_4 ( .A(N436), .Z(out_o[0]) );
endmodule


module mux ( .data_i({\data_i[31][31] , \data_i[31][30] , \data_i[31][29] , 
        \data_i[31][28] , \data_i[31][27] , \data_i[31][26] , \data_i[31][25] , 
        \data_i[31][24] , \data_i[31][23] , \data_i[31][22] , \data_i[31][21] , 
        \data_i[31][20] , \data_i[31][19] , \data_i[31][18] , \data_i[31][17] , 
        \data_i[31][16] , \data_i[31][15] , \data_i[31][14] , \data_i[31][13] , 
        \data_i[31][12] , \data_i[31][11] , \data_i[31][10] , \data_i[31][9] , 
        \data_i[31][8] , \data_i[31][7] , \data_i[31][6] , \data_i[31][5] , 
        \data_i[31][4] , \data_i[31][3] , \data_i[31][2] , \data_i[31][1] , 
        \data_i[31][0] , \data_i[30][31] , \data_i[30][30] , \data_i[30][29] , 
        \data_i[30][28] , \data_i[30][27] , \data_i[30][26] , \data_i[30][25] , 
        \data_i[30][24] , \data_i[30][23] , \data_i[30][22] , \data_i[30][21] , 
        \data_i[30][20] , \data_i[30][19] , \data_i[30][18] , \data_i[30][17] , 
        \data_i[30][16] , \data_i[30][15] , \data_i[30][14] , \data_i[30][13] , 
        \data_i[30][12] , \data_i[30][11] , \data_i[30][10] , \data_i[30][9] , 
        \data_i[30][8] , \data_i[30][7] , \data_i[30][6] , \data_i[30][5] , 
        \data_i[30][4] , \data_i[30][3] , \data_i[30][2] , \data_i[30][1] , 
        \data_i[30][0] , \data_i[29][31] , \data_i[29][30] , \data_i[29][29] , 
        \data_i[29][28] , \data_i[29][27] , \data_i[29][26] , \data_i[29][25] , 
        \data_i[29][24] , \data_i[29][23] , \data_i[29][22] , \data_i[29][21] , 
        \data_i[29][20] , \data_i[29][19] , \data_i[29][18] , \data_i[29][17] , 
        \data_i[29][16] , \data_i[29][15] , \data_i[29][14] , \data_i[29][13] , 
        \data_i[29][12] , \data_i[29][11] , \data_i[29][10] , \data_i[29][9] , 
        \data_i[29][8] , \data_i[29][7] , \data_i[29][6] , \data_i[29][5] , 
        \data_i[29][4] , \data_i[29][3] , \data_i[29][2] , \data_i[29][1] , 
        \data_i[29][0] , \data_i[28][31] , \data_i[28][30] , \data_i[28][29] , 
        \data_i[28][28] , \data_i[28][27] , \data_i[28][26] , \data_i[28][25] , 
        \data_i[28][24] , \data_i[28][23] , \data_i[28][22] , \data_i[28][21] , 
        \data_i[28][20] , \data_i[28][19] , \data_i[28][18] , \data_i[28][17] , 
        \data_i[28][16] , \data_i[28][15] , \data_i[28][14] , \data_i[28][13] , 
        \data_i[28][12] , \data_i[28][11] , \data_i[28][10] , \data_i[28][9] , 
        \data_i[28][8] , \data_i[28][7] , \data_i[28][6] , \data_i[28][5] , 
        \data_i[28][4] , \data_i[28][3] , \data_i[28][2] , \data_i[28][1] , 
        \data_i[28][0] , \data_i[27][31] , \data_i[27][30] , \data_i[27][29] , 
        \data_i[27][28] , \data_i[27][27] , \data_i[27][26] , \data_i[27][25] , 
        \data_i[27][24] , \data_i[27][23] , \data_i[27][22] , \data_i[27][21] , 
        \data_i[27][20] , \data_i[27][19] , \data_i[27][18] , \data_i[27][17] , 
        \data_i[27][16] , \data_i[27][15] , \data_i[27][14] , \data_i[27][13] , 
        \data_i[27][12] , \data_i[27][11] , \data_i[27][10] , \data_i[27][9] , 
        \data_i[27][8] , \data_i[27][7] , \data_i[27][6] , \data_i[27][5] , 
        \data_i[27][4] , \data_i[27][3] , \data_i[27][2] , \data_i[27][1] , 
        \data_i[27][0] , \data_i[26][31] , \data_i[26][30] , \data_i[26][29] , 
        \data_i[26][28] , \data_i[26][27] , \data_i[26][26] , \data_i[26][25] , 
        \data_i[26][24] , \data_i[26][23] , \data_i[26][22] , \data_i[26][21] , 
        \data_i[26][20] , \data_i[26][19] , \data_i[26][18] , \data_i[26][17] , 
        \data_i[26][16] , \data_i[26][15] , \data_i[26][14] , \data_i[26][13] , 
        \data_i[26][12] , \data_i[26][11] , \data_i[26][10] , \data_i[26][9] , 
        \data_i[26][8] , \data_i[26][7] , \data_i[26][6] , \data_i[26][5] , 
        \data_i[26][4] , \data_i[26][3] , \data_i[26][2] , \data_i[26][1] , 
        \data_i[26][0] , \data_i[25][31] , \data_i[25][30] , \data_i[25][29] , 
        \data_i[25][28] , \data_i[25][27] , \data_i[25][26] , \data_i[25][25] , 
        \data_i[25][24] , \data_i[25][23] , \data_i[25][22] , \data_i[25][21] , 
        \data_i[25][20] , \data_i[25][19] , \data_i[25][18] , \data_i[25][17] , 
        \data_i[25][16] , \data_i[25][15] , \data_i[25][14] , \data_i[25][13] , 
        \data_i[25][12] , \data_i[25][11] , \data_i[25][10] , \data_i[25][9] , 
        \data_i[25][8] , \data_i[25][7] , \data_i[25][6] , \data_i[25][5] , 
        \data_i[25][4] , \data_i[25][3] , \data_i[25][2] , \data_i[25][1] , 
        \data_i[25][0] , \data_i[24][31] , \data_i[24][30] , \data_i[24][29] , 
        \data_i[24][28] , \data_i[24][27] , \data_i[24][26] , \data_i[24][25] , 
        \data_i[24][24] , \data_i[24][23] , \data_i[24][22] , \data_i[24][21] , 
        \data_i[24][20] , \data_i[24][19] , \data_i[24][18] , \data_i[24][17] , 
        \data_i[24][16] , \data_i[24][15] , \data_i[24][14] , \data_i[24][13] , 
        \data_i[24][12] , \data_i[24][11] , \data_i[24][10] , \data_i[24][9] , 
        \data_i[24][8] , \data_i[24][7] , \data_i[24][6] , \data_i[24][5] , 
        \data_i[24][4] , \data_i[24][3] , \data_i[24][2] , \data_i[24][1] , 
        \data_i[24][0] , \data_i[23][31] , \data_i[23][30] , \data_i[23][29] , 
        \data_i[23][28] , \data_i[23][27] , \data_i[23][26] , \data_i[23][25] , 
        \data_i[23][24] , \data_i[23][23] , \data_i[23][22] , \data_i[23][21] , 
        \data_i[23][20] , \data_i[23][19] , \data_i[23][18] , \data_i[23][17] , 
        \data_i[23][16] , \data_i[23][15] , \data_i[23][14] , \data_i[23][13] , 
        \data_i[23][12] , \data_i[23][11] , \data_i[23][10] , \data_i[23][9] , 
        \data_i[23][8] , \data_i[23][7] , \data_i[23][6] , \data_i[23][5] , 
        \data_i[23][4] , \data_i[23][3] , \data_i[23][2] , \data_i[23][1] , 
        \data_i[23][0] , \data_i[22][31] , \data_i[22][30] , \data_i[22][29] , 
        \data_i[22][28] , \data_i[22][27] , \data_i[22][26] , \data_i[22][25] , 
        \data_i[22][24] , \data_i[22][23] , \data_i[22][22] , \data_i[22][21] , 
        \data_i[22][20] , \data_i[22][19] , \data_i[22][18] , \data_i[22][17] , 
        \data_i[22][16] , \data_i[22][15] , \data_i[22][14] , \data_i[22][13] , 
        \data_i[22][12] , \data_i[22][11] , \data_i[22][10] , \data_i[22][9] , 
        \data_i[22][8] , \data_i[22][7] , \data_i[22][6] , \data_i[22][5] , 
        \data_i[22][4] , \data_i[22][3] , \data_i[22][2] , \data_i[22][1] , 
        \data_i[22][0] , \data_i[21][31] , \data_i[21][30] , \data_i[21][29] , 
        \data_i[21][28] , \data_i[21][27] , \data_i[21][26] , \data_i[21][25] , 
        \data_i[21][24] , \data_i[21][23] , \data_i[21][22] , \data_i[21][21] , 
        \data_i[21][20] , \data_i[21][19] , \data_i[21][18] , \data_i[21][17] , 
        \data_i[21][16] , \data_i[21][15] , \data_i[21][14] , \data_i[21][13] , 
        \data_i[21][12] , \data_i[21][11] , \data_i[21][10] , \data_i[21][9] , 
        \data_i[21][8] , \data_i[21][7] , \data_i[21][6] , \data_i[21][5] , 
        \data_i[21][4] , \data_i[21][3] , \data_i[21][2] , \data_i[21][1] , 
        \data_i[21][0] , \data_i[20][31] , \data_i[20][30] , \data_i[20][29] , 
        \data_i[20][28] , \data_i[20][27] , \data_i[20][26] , \data_i[20][25] , 
        \data_i[20][24] , \data_i[20][23] , \data_i[20][22] , \data_i[20][21] , 
        \data_i[20][20] , \data_i[20][19] , \data_i[20][18] , \data_i[20][17] , 
        \data_i[20][16] , \data_i[20][15] , \data_i[20][14] , \data_i[20][13] , 
        \data_i[20][12] , \data_i[20][11] , \data_i[20][10] , \data_i[20][9] , 
        \data_i[20][8] , \data_i[20][7] , \data_i[20][6] , \data_i[20][5] , 
        \data_i[20][4] , \data_i[20][3] , \data_i[20][2] , \data_i[20][1] , 
        \data_i[20][0] , \data_i[19][31] , \data_i[19][30] , \data_i[19][29] , 
        \data_i[19][28] , \data_i[19][27] , \data_i[19][26] , \data_i[19][25] , 
        \data_i[19][24] , \data_i[19][23] , \data_i[19][22] , \data_i[19][21] , 
        \data_i[19][20] , \data_i[19][19] , \data_i[19][18] , \data_i[19][17] , 
        \data_i[19][16] , \data_i[19][15] , \data_i[19][14] , \data_i[19][13] , 
        \data_i[19][12] , \data_i[19][11] , \data_i[19][10] , \data_i[19][9] , 
        \data_i[19][8] , \data_i[19][7] , \data_i[19][6] , \data_i[19][5] , 
        \data_i[19][4] , \data_i[19][3] , \data_i[19][2] , \data_i[19][1] , 
        \data_i[19][0] , \data_i[18][31] , \data_i[18][30] , \data_i[18][29] , 
        \data_i[18][28] , \data_i[18][27] , \data_i[18][26] , \data_i[18][25] , 
        \data_i[18][24] , \data_i[18][23] , \data_i[18][22] , \data_i[18][21] , 
        \data_i[18][20] , \data_i[18][19] , \data_i[18][18] , \data_i[18][17] , 
        \data_i[18][16] , \data_i[18][15] , \data_i[18][14] , \data_i[18][13] , 
        \data_i[18][12] , \data_i[18][11] , \data_i[18][10] , \data_i[18][9] , 
        \data_i[18][8] , \data_i[18][7] , \data_i[18][6] , \data_i[18][5] , 
        \data_i[18][4] , \data_i[18][3] , \data_i[18][2] , \data_i[18][1] , 
        \data_i[18][0] , \data_i[17][31] , \data_i[17][30] , \data_i[17][29] , 
        \data_i[17][28] , \data_i[17][27] , \data_i[17][26] , \data_i[17][25] , 
        \data_i[17][24] , \data_i[17][23] , \data_i[17][22] , \data_i[17][21] , 
        \data_i[17][20] , \data_i[17][19] , \data_i[17][18] , \data_i[17][17] , 
        \data_i[17][16] , \data_i[17][15] , \data_i[17][14] , \data_i[17][13] , 
        \data_i[17][12] , \data_i[17][11] , \data_i[17][10] , \data_i[17][9] , 
        \data_i[17][8] , \data_i[17][7] , \data_i[17][6] , \data_i[17][5] , 
        \data_i[17][4] , \data_i[17][3] , \data_i[17][2] , \data_i[17][1] , 
        \data_i[17][0] , \data_i[16][31] , \data_i[16][30] , \data_i[16][29] , 
        \data_i[16][28] , \data_i[16][27] , \data_i[16][26] , \data_i[16][25] , 
        \data_i[16][24] , \data_i[16][23] , \data_i[16][22] , \data_i[16][21] , 
        \data_i[16][20] , \data_i[16][19] , \data_i[16][18] , \data_i[16][17] , 
        \data_i[16][16] , \data_i[16][15] , \data_i[16][14] , \data_i[16][13] , 
        \data_i[16][12] , \data_i[16][11] , \data_i[16][10] , \data_i[16][9] , 
        \data_i[16][8] , \data_i[16][7] , \data_i[16][6] , \data_i[16][5] , 
        \data_i[16][4] , \data_i[16][3] , \data_i[16][2] , \data_i[16][1] , 
        \data_i[16][0] , \data_i[15][31] , \data_i[15][30] , \data_i[15][29] , 
        \data_i[15][28] , \data_i[15][27] , \data_i[15][26] , \data_i[15][25] , 
        \data_i[15][24] , \data_i[15][23] , \data_i[15][22] , \data_i[15][21] , 
        \data_i[15][20] , \data_i[15][19] , \data_i[15][18] , \data_i[15][17] , 
        \data_i[15][16] , \data_i[15][15] , \data_i[15][14] , \data_i[15][13] , 
        \data_i[15][12] , \data_i[15][11] , \data_i[15][10] , \data_i[15][9] , 
        \data_i[15][8] , \data_i[15][7] , \data_i[15][6] , \data_i[15][5] , 
        \data_i[15][4] , \data_i[15][3] , \data_i[15][2] , \data_i[15][1] , 
        \data_i[15][0] , \data_i[14][31] , \data_i[14][30] , \data_i[14][29] , 
        \data_i[14][28] , \data_i[14][27] , \data_i[14][26] , \data_i[14][25] , 
        \data_i[14][24] , \data_i[14][23] , \data_i[14][22] , \data_i[14][21] , 
        \data_i[14][20] , \data_i[14][19] , \data_i[14][18] , \data_i[14][17] , 
        \data_i[14][16] , \data_i[14][15] , \data_i[14][14] , \data_i[14][13] , 
        \data_i[14][12] , \data_i[14][11] , \data_i[14][10] , \data_i[14][9] , 
        \data_i[14][8] , \data_i[14][7] , \data_i[14][6] , \data_i[14][5] , 
        \data_i[14][4] , \data_i[14][3] , \data_i[14][2] , \data_i[14][1] , 
        \data_i[14][0] , \data_i[13][31] , \data_i[13][30] , \data_i[13][29] , 
        \data_i[13][28] , \data_i[13][27] , \data_i[13][26] , \data_i[13][25] , 
        \data_i[13][24] , \data_i[13][23] , \data_i[13][22] , \data_i[13][21] , 
        \data_i[13][20] , \data_i[13][19] , \data_i[13][18] , \data_i[13][17] , 
        \data_i[13][16] , \data_i[13][15] , \data_i[13][14] , \data_i[13][13] , 
        \data_i[13][12] , \data_i[13][11] , \data_i[13][10] , \data_i[13][9] , 
        \data_i[13][8] , \data_i[13][7] , \data_i[13][6] , \data_i[13][5] , 
        \data_i[13][4] , \data_i[13][3] , \data_i[13][2] , \data_i[13][1] , 
        \data_i[13][0] , \data_i[12][31] , \data_i[12][30] , \data_i[12][29] , 
        \data_i[12][28] , \data_i[12][27] , \data_i[12][26] , \data_i[12][25] , 
        \data_i[12][24] , \data_i[12][23] , \data_i[12][22] , \data_i[12][21] , 
        \data_i[12][20] , \data_i[12][19] , \data_i[12][18] , \data_i[12][17] , 
        \data_i[12][16] , \data_i[12][15] , \data_i[12][14] , \data_i[12][13] , 
        \data_i[12][12] , \data_i[12][11] , \data_i[12][10] , \data_i[12][9] , 
        \data_i[12][8] , \data_i[12][7] , \data_i[12][6] , \data_i[12][5] , 
        \data_i[12][4] , \data_i[12][3] , \data_i[12][2] , \data_i[12][1] , 
        \data_i[12][0] , \data_i[11][31] , \data_i[11][30] , \data_i[11][29] , 
        \data_i[11][28] , \data_i[11][27] , \data_i[11][26] , \data_i[11][25] , 
        \data_i[11][24] , \data_i[11][23] , \data_i[11][22] , \data_i[11][21] , 
        \data_i[11][20] , \data_i[11][19] , \data_i[11][18] , \data_i[11][17] , 
        \data_i[11][16] , \data_i[11][15] , \data_i[11][14] , \data_i[11][13] , 
        \data_i[11][12] , \data_i[11][11] , \data_i[11][10] , \data_i[11][9] , 
        \data_i[11][8] , \data_i[11][7] , \data_i[11][6] , \data_i[11][5] , 
        \data_i[11][4] , \data_i[11][3] , \data_i[11][2] , \data_i[11][1] , 
        \data_i[11][0] , \data_i[10][31] , \data_i[10][30] , \data_i[10][29] , 
        \data_i[10][28] , \data_i[10][27] , \data_i[10][26] , \data_i[10][25] , 
        \data_i[10][24] , \data_i[10][23] , \data_i[10][22] , \data_i[10][21] , 
        \data_i[10][20] , \data_i[10][19] , \data_i[10][18] , \data_i[10][17] , 
        \data_i[10][16] , \data_i[10][15] , \data_i[10][14] , \data_i[10][13] , 
        \data_i[10][12] , \data_i[10][11] , \data_i[10][10] , \data_i[10][9] , 
        \data_i[10][8] , \data_i[10][7] , \data_i[10][6] , \data_i[10][5] , 
        \data_i[10][4] , \data_i[10][3] , \data_i[10][2] , \data_i[10][1] , 
        \data_i[10][0] , \data_i[9][31] , \data_i[9][30] , \data_i[9][29] , 
        \data_i[9][28] , \data_i[9][27] , \data_i[9][26] , \data_i[9][25] , 
        \data_i[9][24] , \data_i[9][23] , \data_i[9][22] , \data_i[9][21] , 
        \data_i[9][20] , \data_i[9][19] , \data_i[9][18] , \data_i[9][17] , 
        \data_i[9][16] , \data_i[9][15] , \data_i[9][14] , \data_i[9][13] , 
        \data_i[9][12] , \data_i[9][11] , \data_i[9][10] , \data_i[9][9] , 
        \data_i[9][8] , \data_i[9][7] , \data_i[9][6] , \data_i[9][5] , 
        \data_i[9][4] , \data_i[9][3] , \data_i[9][2] , \data_i[9][1] , 
        \data_i[9][0] , \data_i[8][31] , \data_i[8][30] , \data_i[8][29] , 
        \data_i[8][28] , \data_i[8][27] , \data_i[8][26] , \data_i[8][25] , 
        \data_i[8][24] , \data_i[8][23] , \data_i[8][22] , \data_i[8][21] , 
        \data_i[8][20] , \data_i[8][19] , \data_i[8][18] , \data_i[8][17] , 
        \data_i[8][16] , \data_i[8][15] , \data_i[8][14] , \data_i[8][13] , 
        \data_i[8][12] , \data_i[8][11] , \data_i[8][10] , \data_i[8][9] , 
        \data_i[8][8] , \data_i[8][7] , \data_i[8][6] , \data_i[8][5] , 
        \data_i[8][4] , \data_i[8][3] , \data_i[8][2] , \data_i[8][1] , 
        \data_i[8][0] , \data_i[7][31] , \data_i[7][30] , \data_i[7][29] , 
        \data_i[7][28] , \data_i[7][27] , \data_i[7][26] , \data_i[7][25] , 
        \data_i[7][24] , \data_i[7][23] , \data_i[7][22] , \data_i[7][21] , 
        \data_i[7][20] , \data_i[7][19] , \data_i[7][18] , \data_i[7][17] , 
        \data_i[7][16] , \data_i[7][15] , \data_i[7][14] , \data_i[7][13] , 
        \data_i[7][12] , \data_i[7][11] , \data_i[7][10] , \data_i[7][9] , 
        \data_i[7][8] , \data_i[7][7] , \data_i[7][6] , \data_i[7][5] , 
        \data_i[7][4] , \data_i[7][3] , \data_i[7][2] , \data_i[7][1] , 
        \data_i[7][0] , \data_i[6][31] , \data_i[6][30] , \data_i[6][29] , 
        \data_i[6][28] , \data_i[6][27] , \data_i[6][26] , \data_i[6][25] , 
        \data_i[6][24] , \data_i[6][23] , \data_i[6][22] , \data_i[6][21] , 
        \data_i[6][20] , \data_i[6][19] , \data_i[6][18] , \data_i[6][17] , 
        \data_i[6][16] , \data_i[6][15] , \data_i[6][14] , \data_i[6][13] , 
        \data_i[6][12] , \data_i[6][11] , \data_i[6][10] , \data_i[6][9] , 
        \data_i[6][8] , \data_i[6][7] , \data_i[6][6] , \data_i[6][5] , 
        \data_i[6][4] , \data_i[6][3] , \data_i[6][2] , \data_i[6][1] , 
        \data_i[6][0] , \data_i[5][31] , \data_i[5][30] , \data_i[5][29] , 
        \data_i[5][28] , \data_i[5][27] , \data_i[5][26] , \data_i[5][25] , 
        \data_i[5][24] , \data_i[5][23] , \data_i[5][22] , \data_i[5][21] , 
        \data_i[5][20] , \data_i[5][19] , \data_i[5][18] , \data_i[5][17] , 
        \data_i[5][16] , \data_i[5][15] , \data_i[5][14] , \data_i[5][13] , 
        \data_i[5][12] , \data_i[5][11] , \data_i[5][10] , \data_i[5][9] , 
        \data_i[5][8] , \data_i[5][7] , \data_i[5][6] , \data_i[5][5] , 
        \data_i[5][4] , \data_i[5][3] , \data_i[5][2] , \data_i[5][1] , 
        \data_i[5][0] , \data_i[4][31] , \data_i[4][30] , \data_i[4][29] , 
        \data_i[4][28] , \data_i[4][27] , \data_i[4][26] , \data_i[4][25] , 
        \data_i[4][24] , \data_i[4][23] , \data_i[4][22] , \data_i[4][21] , 
        \data_i[4][20] , \data_i[4][19] , \data_i[4][18] , \data_i[4][17] , 
        \data_i[4][16] , \data_i[4][15] , \data_i[4][14] , \data_i[4][13] , 
        \data_i[4][12] , \data_i[4][11] , \data_i[4][10] , \data_i[4][9] , 
        \data_i[4][8] , \data_i[4][7] , \data_i[4][6] , \data_i[4][5] , 
        \data_i[4][4] , \data_i[4][3] , \data_i[4][2] , \data_i[4][1] , 
        \data_i[4][0] , \data_i[3][31] , \data_i[3][30] , \data_i[3][29] , 
        \data_i[3][28] , \data_i[3][27] , \data_i[3][26] , \data_i[3][25] , 
        \data_i[3][24] , \data_i[3][23] , \data_i[3][22] , \data_i[3][21] , 
        \data_i[3][20] , \data_i[3][19] , \data_i[3][18] , \data_i[3][17] , 
        \data_i[3][16] , \data_i[3][15] , \data_i[3][14] , \data_i[3][13] , 
        \data_i[3][12] , \data_i[3][11] , \data_i[3][10] , \data_i[3][9] , 
        \data_i[3][8] , \data_i[3][7] , \data_i[3][6] , \data_i[3][5] , 
        \data_i[3][4] , \data_i[3][3] , \data_i[3][2] , \data_i[3][1] , 
        \data_i[3][0] , \data_i[2][31] , \data_i[2][30] , \data_i[2][29] , 
        \data_i[2][28] , \data_i[2][27] , \data_i[2][26] , \data_i[2][25] , 
        \data_i[2][24] , \data_i[2][23] , \data_i[2][22] , \data_i[2][21] , 
        \data_i[2][20] , \data_i[2][19] , \data_i[2][18] , \data_i[2][17] , 
        \data_i[2][16] , \data_i[2][15] , \data_i[2][14] , \data_i[2][13] , 
        \data_i[2][12] , \data_i[2][11] , \data_i[2][10] , \data_i[2][9] , 
        \data_i[2][8] , \data_i[2][7] , \data_i[2][6] , \data_i[2][5] , 
        \data_i[2][4] , \data_i[2][3] , \data_i[2][2] , \data_i[2][1] , 
        \data_i[2][0] , \data_i[1][31] , \data_i[1][30] , \data_i[1][29] , 
        \data_i[1][28] , \data_i[1][27] , \data_i[1][26] , \data_i[1][25] , 
        \data_i[1][24] , \data_i[1][23] , \data_i[1][22] , \data_i[1][21] , 
        \data_i[1][20] , \data_i[1][19] , \data_i[1][18] , \data_i[1][17] , 
        \data_i[1][16] , \data_i[1][15] , \data_i[1][14] , \data_i[1][13] , 
        \data_i[1][12] , \data_i[1][11] , \data_i[1][10] , \data_i[1][9] , 
        \data_i[1][8] , \data_i[1][7] , \data_i[1][6] , \data_i[1][5] , 
        \data_i[1][4] , \data_i[1][3] , \data_i[1][2] , \data_i[1][1] , 
        \data_i[1][0] , \data_i[0][31] , \data_i[0][30] , \data_i[0][29] , 
        \data_i[0][28] , \data_i[0][27] , \data_i[0][26] , \data_i[0][25] , 
        \data_i[0][24] , \data_i[0][23] , \data_i[0][22] , \data_i[0][21] , 
        \data_i[0][20] , \data_i[0][19] , \data_i[0][18] , \data_i[0][17] , 
        \data_i[0][16] , \data_i[0][15] , \data_i[0][14] , \data_i[0][13] , 
        \data_i[0][12] , \data_i[0][11] , \data_i[0][10] , \data_i[0][9] , 
        \data_i[0][8] , \data_i[0][7] , \data_i[0][6] , \data_i[0][5] , 
        \data_i[0][4] , \data_i[0][3] , \data_i[0][2] , \data_i[0][1] , 
        \data_i[0][0] }), select_i, data_o );
  input [4:0] select_i;
  output [31:0] data_o;
  input \data_i[31][31] , \data_i[31][30] , \data_i[31][29] , \data_i[31][28] ,
         \data_i[31][27] , \data_i[31][26] , \data_i[31][25] ,
         \data_i[31][24] , \data_i[31][23] , \data_i[31][22] ,
         \data_i[31][21] , \data_i[31][20] , \data_i[31][19] ,
         \data_i[31][18] , \data_i[31][17] , \data_i[31][16] ,
         \data_i[31][15] , \data_i[31][14] , \data_i[31][13] ,
         \data_i[31][12] , \data_i[31][11] , \data_i[31][10] , \data_i[31][9] ,
         \data_i[31][8] , \data_i[31][7] , \data_i[31][6] , \data_i[31][5] ,
         \data_i[31][4] , \data_i[31][3] , \data_i[31][2] , \data_i[31][1] ,
         \data_i[31][0] , \data_i[30][31] , \data_i[30][30] , \data_i[30][29] ,
         \data_i[30][28] , \data_i[30][27] , \data_i[30][26] ,
         \data_i[30][25] , \data_i[30][24] , \data_i[30][23] ,
         \data_i[30][22] , \data_i[30][21] , \data_i[30][20] ,
         \data_i[30][19] , \data_i[30][18] , \data_i[30][17] ,
         \data_i[30][16] , \data_i[30][15] , \data_i[30][14] ,
         \data_i[30][13] , \data_i[30][12] , \data_i[30][11] ,
         \data_i[30][10] , \data_i[30][9] , \data_i[30][8] , \data_i[30][7] ,
         \data_i[30][6] , \data_i[30][5] , \data_i[30][4] , \data_i[30][3] ,
         \data_i[30][2] , \data_i[30][1] , \data_i[30][0] , \data_i[29][31] ,
         \data_i[29][30] , \data_i[29][29] , \data_i[29][28] ,
         \data_i[29][27] , \data_i[29][26] , \data_i[29][25] ,
         \data_i[29][24] , \data_i[29][23] , \data_i[29][22] ,
         \data_i[29][21] , \data_i[29][20] , \data_i[29][19] ,
         \data_i[29][18] , \data_i[29][17] , \data_i[29][16] ,
         \data_i[29][15] , \data_i[29][14] , \data_i[29][13] ,
         \data_i[29][12] , \data_i[29][11] , \data_i[29][10] , \data_i[29][9] ,
         \data_i[29][8] , \data_i[29][7] , \data_i[29][6] , \data_i[29][5] ,
         \data_i[29][4] , \data_i[29][3] , \data_i[29][2] , \data_i[29][1] ,
         \data_i[29][0] , \data_i[28][31] , \data_i[28][30] , \data_i[28][29] ,
         \data_i[28][28] , \data_i[28][27] , \data_i[28][26] ,
         \data_i[28][25] , \data_i[28][24] , \data_i[28][23] ,
         \data_i[28][22] , \data_i[28][21] , \data_i[28][20] ,
         \data_i[28][19] , \data_i[28][18] , \data_i[28][17] ,
         \data_i[28][16] , \data_i[28][15] , \data_i[28][14] ,
         \data_i[28][13] , \data_i[28][12] , \data_i[28][11] ,
         \data_i[28][10] , \data_i[28][9] , \data_i[28][8] , \data_i[28][7] ,
         \data_i[28][6] , \data_i[28][5] , \data_i[28][4] , \data_i[28][3] ,
         \data_i[28][2] , \data_i[28][1] , \data_i[28][0] , \data_i[27][31] ,
         \data_i[27][30] , \data_i[27][29] , \data_i[27][28] ,
         \data_i[27][27] , \data_i[27][26] , \data_i[27][25] ,
         \data_i[27][24] , \data_i[27][23] , \data_i[27][22] ,
         \data_i[27][21] , \data_i[27][20] , \data_i[27][19] ,
         \data_i[27][18] , \data_i[27][17] , \data_i[27][16] ,
         \data_i[27][15] , \data_i[27][14] , \data_i[27][13] ,
         \data_i[27][12] , \data_i[27][11] , \data_i[27][10] , \data_i[27][9] ,
         \data_i[27][8] , \data_i[27][7] , \data_i[27][6] , \data_i[27][5] ,
         \data_i[27][4] , \data_i[27][3] , \data_i[27][2] , \data_i[27][1] ,
         \data_i[27][0] , \data_i[26][31] , \data_i[26][30] , \data_i[26][29] ,
         \data_i[26][28] , \data_i[26][27] , \data_i[26][26] ,
         \data_i[26][25] , \data_i[26][24] , \data_i[26][23] ,
         \data_i[26][22] , \data_i[26][21] , \data_i[26][20] ,
         \data_i[26][19] , \data_i[26][18] , \data_i[26][17] ,
         \data_i[26][16] , \data_i[26][15] , \data_i[26][14] ,
         \data_i[26][13] , \data_i[26][12] , \data_i[26][11] ,
         \data_i[26][10] , \data_i[26][9] , \data_i[26][8] , \data_i[26][7] ,
         \data_i[26][6] , \data_i[26][5] , \data_i[26][4] , \data_i[26][3] ,
         \data_i[26][2] , \data_i[26][1] , \data_i[26][0] , \data_i[25][31] ,
         \data_i[25][30] , \data_i[25][29] , \data_i[25][28] ,
         \data_i[25][27] , \data_i[25][26] , \data_i[25][25] ,
         \data_i[25][24] , \data_i[25][23] , \data_i[25][22] ,
         \data_i[25][21] , \data_i[25][20] , \data_i[25][19] ,
         \data_i[25][18] , \data_i[25][17] , \data_i[25][16] ,
         \data_i[25][15] , \data_i[25][14] , \data_i[25][13] ,
         \data_i[25][12] , \data_i[25][11] , \data_i[25][10] , \data_i[25][9] ,
         \data_i[25][8] , \data_i[25][7] , \data_i[25][6] , \data_i[25][5] ,
         \data_i[25][4] , \data_i[25][3] , \data_i[25][2] , \data_i[25][1] ,
         \data_i[25][0] , \data_i[24][31] , \data_i[24][30] , \data_i[24][29] ,
         \data_i[24][28] , \data_i[24][27] , \data_i[24][26] ,
         \data_i[24][25] , \data_i[24][24] , \data_i[24][23] ,
         \data_i[24][22] , \data_i[24][21] , \data_i[24][20] ,
         \data_i[24][19] , \data_i[24][18] , \data_i[24][17] ,
         \data_i[24][16] , \data_i[24][15] , \data_i[24][14] ,
         \data_i[24][13] , \data_i[24][12] , \data_i[24][11] ,
         \data_i[24][10] , \data_i[24][9] , \data_i[24][8] , \data_i[24][7] ,
         \data_i[24][6] , \data_i[24][5] , \data_i[24][4] , \data_i[24][3] ,
         \data_i[24][2] , \data_i[24][1] , \data_i[24][0] , \data_i[23][31] ,
         \data_i[23][30] , \data_i[23][29] , \data_i[23][28] ,
         \data_i[23][27] , \data_i[23][26] , \data_i[23][25] ,
         \data_i[23][24] , \data_i[23][23] , \data_i[23][22] ,
         \data_i[23][21] , \data_i[23][20] , \data_i[23][19] ,
         \data_i[23][18] , \data_i[23][17] , \data_i[23][16] ,
         \data_i[23][15] , \data_i[23][14] , \data_i[23][13] ,
         \data_i[23][12] , \data_i[23][11] , \data_i[23][10] , \data_i[23][9] ,
         \data_i[23][8] , \data_i[23][7] , \data_i[23][6] , \data_i[23][5] ,
         \data_i[23][4] , \data_i[23][3] , \data_i[23][2] , \data_i[23][1] ,
         \data_i[23][0] , \data_i[22][31] , \data_i[22][30] , \data_i[22][29] ,
         \data_i[22][28] , \data_i[22][27] , \data_i[22][26] ,
         \data_i[22][25] , \data_i[22][24] , \data_i[22][23] ,
         \data_i[22][22] , \data_i[22][21] , \data_i[22][20] ,
         \data_i[22][19] , \data_i[22][18] , \data_i[22][17] ,
         \data_i[22][16] , \data_i[22][15] , \data_i[22][14] ,
         \data_i[22][13] , \data_i[22][12] , \data_i[22][11] ,
         \data_i[22][10] , \data_i[22][9] , \data_i[22][8] , \data_i[22][7] ,
         \data_i[22][6] , \data_i[22][5] , \data_i[22][4] , \data_i[22][3] ,
         \data_i[22][2] , \data_i[22][1] , \data_i[22][0] , \data_i[21][31] ,
         \data_i[21][30] , \data_i[21][29] , \data_i[21][28] ,
         \data_i[21][27] , \data_i[21][26] , \data_i[21][25] ,
         \data_i[21][24] , \data_i[21][23] , \data_i[21][22] ,
         \data_i[21][21] , \data_i[21][20] , \data_i[21][19] ,
         \data_i[21][18] , \data_i[21][17] , \data_i[21][16] ,
         \data_i[21][15] , \data_i[21][14] , \data_i[21][13] ,
         \data_i[21][12] , \data_i[21][11] , \data_i[21][10] , \data_i[21][9] ,
         \data_i[21][8] , \data_i[21][7] , \data_i[21][6] , \data_i[21][5] ,
         \data_i[21][4] , \data_i[21][3] , \data_i[21][2] , \data_i[21][1] ,
         \data_i[21][0] , \data_i[20][31] , \data_i[20][30] , \data_i[20][29] ,
         \data_i[20][28] , \data_i[20][27] , \data_i[20][26] ,
         \data_i[20][25] , \data_i[20][24] , \data_i[20][23] ,
         \data_i[20][22] , \data_i[20][21] , \data_i[20][20] ,
         \data_i[20][19] , \data_i[20][18] , \data_i[20][17] ,
         \data_i[20][16] , \data_i[20][15] , \data_i[20][14] ,
         \data_i[20][13] , \data_i[20][12] , \data_i[20][11] ,
         \data_i[20][10] , \data_i[20][9] , \data_i[20][8] , \data_i[20][7] ,
         \data_i[20][6] , \data_i[20][5] , \data_i[20][4] , \data_i[20][3] ,
         \data_i[20][2] , \data_i[20][1] , \data_i[20][0] , \data_i[19][31] ,
         \data_i[19][30] , \data_i[19][29] , \data_i[19][28] ,
         \data_i[19][27] , \data_i[19][26] , \data_i[19][25] ,
         \data_i[19][24] , \data_i[19][23] , \data_i[19][22] ,
         \data_i[19][21] , \data_i[19][20] , \data_i[19][19] ,
         \data_i[19][18] , \data_i[19][17] , \data_i[19][16] ,
         \data_i[19][15] , \data_i[19][14] , \data_i[19][13] ,
         \data_i[19][12] , \data_i[19][11] , \data_i[19][10] , \data_i[19][9] ,
         \data_i[19][8] , \data_i[19][7] , \data_i[19][6] , \data_i[19][5] ,
         \data_i[19][4] , \data_i[19][3] , \data_i[19][2] , \data_i[19][1] ,
         \data_i[19][0] , \data_i[18][31] , \data_i[18][30] , \data_i[18][29] ,
         \data_i[18][28] , \data_i[18][27] , \data_i[18][26] ,
         \data_i[18][25] , \data_i[18][24] , \data_i[18][23] ,
         \data_i[18][22] , \data_i[18][21] , \data_i[18][20] ,
         \data_i[18][19] , \data_i[18][18] , \data_i[18][17] ,
         \data_i[18][16] , \data_i[18][15] , \data_i[18][14] ,
         \data_i[18][13] , \data_i[18][12] , \data_i[18][11] ,
         \data_i[18][10] , \data_i[18][9] , \data_i[18][8] , \data_i[18][7] ,
         \data_i[18][6] , \data_i[18][5] , \data_i[18][4] , \data_i[18][3] ,
         \data_i[18][2] , \data_i[18][1] , \data_i[18][0] , \data_i[17][31] ,
         \data_i[17][30] , \data_i[17][29] , \data_i[17][28] ,
         \data_i[17][27] , \data_i[17][26] , \data_i[17][25] ,
         \data_i[17][24] , \data_i[17][23] , \data_i[17][22] ,
         \data_i[17][21] , \data_i[17][20] , \data_i[17][19] ,
         \data_i[17][18] , \data_i[17][17] , \data_i[17][16] ,
         \data_i[17][15] , \data_i[17][14] , \data_i[17][13] ,
         \data_i[17][12] , \data_i[17][11] , \data_i[17][10] , \data_i[17][9] ,
         \data_i[17][8] , \data_i[17][7] , \data_i[17][6] , \data_i[17][5] ,
         \data_i[17][4] , \data_i[17][3] , \data_i[17][2] , \data_i[17][1] ,
         \data_i[17][0] , \data_i[16][31] , \data_i[16][30] , \data_i[16][29] ,
         \data_i[16][28] , \data_i[16][27] , \data_i[16][26] ,
         \data_i[16][25] , \data_i[16][24] , \data_i[16][23] ,
         \data_i[16][22] , \data_i[16][21] , \data_i[16][20] ,
         \data_i[16][19] , \data_i[16][18] , \data_i[16][17] ,
         \data_i[16][16] , \data_i[16][15] , \data_i[16][14] ,
         \data_i[16][13] , \data_i[16][12] , \data_i[16][11] ,
         \data_i[16][10] , \data_i[16][9] , \data_i[16][8] , \data_i[16][7] ,
         \data_i[16][6] , \data_i[16][5] , \data_i[16][4] , \data_i[16][3] ,
         \data_i[16][2] , \data_i[16][1] , \data_i[16][0] , \data_i[15][31] ,
         \data_i[15][30] , \data_i[15][29] , \data_i[15][28] ,
         \data_i[15][27] , \data_i[15][26] , \data_i[15][25] ,
         \data_i[15][24] , \data_i[15][23] , \data_i[15][22] ,
         \data_i[15][21] , \data_i[15][20] , \data_i[15][19] ,
         \data_i[15][18] , \data_i[15][17] , \data_i[15][16] ,
         \data_i[15][15] , \data_i[15][14] , \data_i[15][13] ,
         \data_i[15][12] , \data_i[15][11] , \data_i[15][10] , \data_i[15][9] ,
         \data_i[15][8] , \data_i[15][7] , \data_i[15][6] , \data_i[15][5] ,
         \data_i[15][4] , \data_i[15][3] , \data_i[15][2] , \data_i[15][1] ,
         \data_i[15][0] , \data_i[14][31] , \data_i[14][30] , \data_i[14][29] ,
         \data_i[14][28] , \data_i[14][27] , \data_i[14][26] ,
         \data_i[14][25] , \data_i[14][24] , \data_i[14][23] ,
         \data_i[14][22] , \data_i[14][21] , \data_i[14][20] ,
         \data_i[14][19] , \data_i[14][18] , \data_i[14][17] ,
         \data_i[14][16] , \data_i[14][15] , \data_i[14][14] ,
         \data_i[14][13] , \data_i[14][12] , \data_i[14][11] ,
         \data_i[14][10] , \data_i[14][9] , \data_i[14][8] , \data_i[14][7] ,
         \data_i[14][6] , \data_i[14][5] , \data_i[14][4] , \data_i[14][3] ,
         \data_i[14][2] , \data_i[14][1] , \data_i[14][0] , \data_i[13][31] ,
         \data_i[13][30] , \data_i[13][29] , \data_i[13][28] ,
         \data_i[13][27] , \data_i[13][26] , \data_i[13][25] ,
         \data_i[13][24] , \data_i[13][23] , \data_i[13][22] ,
         \data_i[13][21] , \data_i[13][20] , \data_i[13][19] ,
         \data_i[13][18] , \data_i[13][17] , \data_i[13][16] ,
         \data_i[13][15] , \data_i[13][14] , \data_i[13][13] ,
         \data_i[13][12] , \data_i[13][11] , \data_i[13][10] , \data_i[13][9] ,
         \data_i[13][8] , \data_i[13][7] , \data_i[13][6] , \data_i[13][5] ,
         \data_i[13][4] , \data_i[13][3] , \data_i[13][2] , \data_i[13][1] ,
         \data_i[13][0] , \data_i[12][31] , \data_i[12][30] , \data_i[12][29] ,
         \data_i[12][28] , \data_i[12][27] , \data_i[12][26] ,
         \data_i[12][25] , \data_i[12][24] , \data_i[12][23] ,
         \data_i[12][22] , \data_i[12][21] , \data_i[12][20] ,
         \data_i[12][19] , \data_i[12][18] , \data_i[12][17] ,
         \data_i[12][16] , \data_i[12][15] , \data_i[12][14] ,
         \data_i[12][13] , \data_i[12][12] , \data_i[12][11] ,
         \data_i[12][10] , \data_i[12][9] , \data_i[12][8] , \data_i[12][7] ,
         \data_i[12][6] , \data_i[12][5] , \data_i[12][4] , \data_i[12][3] ,
         \data_i[12][2] , \data_i[12][1] , \data_i[12][0] , \data_i[11][31] ,
         \data_i[11][30] , \data_i[11][29] , \data_i[11][28] ,
         \data_i[11][27] , \data_i[11][26] , \data_i[11][25] ,
         \data_i[11][24] , \data_i[11][23] , \data_i[11][22] ,
         \data_i[11][21] , \data_i[11][20] , \data_i[11][19] ,
         \data_i[11][18] , \data_i[11][17] , \data_i[11][16] ,
         \data_i[11][15] , \data_i[11][14] , \data_i[11][13] ,
         \data_i[11][12] , \data_i[11][11] , \data_i[11][10] , \data_i[11][9] ,
         \data_i[11][8] , \data_i[11][7] , \data_i[11][6] , \data_i[11][5] ,
         \data_i[11][4] , \data_i[11][3] , \data_i[11][2] , \data_i[11][1] ,
         \data_i[11][0] , \data_i[10][31] , \data_i[10][30] , \data_i[10][29] ,
         \data_i[10][28] , \data_i[10][27] , \data_i[10][26] ,
         \data_i[10][25] , \data_i[10][24] , \data_i[10][23] ,
         \data_i[10][22] , \data_i[10][21] , \data_i[10][20] ,
         \data_i[10][19] , \data_i[10][18] , \data_i[10][17] ,
         \data_i[10][16] , \data_i[10][15] , \data_i[10][14] ,
         \data_i[10][13] , \data_i[10][12] , \data_i[10][11] ,
         \data_i[10][10] , \data_i[10][9] , \data_i[10][8] , \data_i[10][7] ,
         \data_i[10][6] , \data_i[10][5] , \data_i[10][4] , \data_i[10][3] ,
         \data_i[10][2] , \data_i[10][1] , \data_i[10][0] , \data_i[9][31] ,
         \data_i[9][30] , \data_i[9][29] , \data_i[9][28] , \data_i[9][27] ,
         \data_i[9][26] , \data_i[9][25] , \data_i[9][24] , \data_i[9][23] ,
         \data_i[9][22] , \data_i[9][21] , \data_i[9][20] , \data_i[9][19] ,
         \data_i[9][18] , \data_i[9][17] , \data_i[9][16] , \data_i[9][15] ,
         \data_i[9][14] , \data_i[9][13] , \data_i[9][12] , \data_i[9][11] ,
         \data_i[9][10] , \data_i[9][9] , \data_i[9][8] , \data_i[9][7] ,
         \data_i[9][6] , \data_i[9][5] , \data_i[9][4] , \data_i[9][3] ,
         \data_i[9][2] , \data_i[9][1] , \data_i[9][0] , \data_i[8][31] ,
         \data_i[8][30] , \data_i[8][29] , \data_i[8][28] , \data_i[8][27] ,
         \data_i[8][26] , \data_i[8][25] , \data_i[8][24] , \data_i[8][23] ,
         \data_i[8][22] , \data_i[8][21] , \data_i[8][20] , \data_i[8][19] ,
         \data_i[8][18] , \data_i[8][17] , \data_i[8][16] , \data_i[8][15] ,
         \data_i[8][14] , \data_i[8][13] , \data_i[8][12] , \data_i[8][11] ,
         \data_i[8][10] , \data_i[8][9] , \data_i[8][8] , \data_i[8][7] ,
         \data_i[8][6] , \data_i[8][5] , \data_i[8][4] , \data_i[8][3] ,
         \data_i[8][2] , \data_i[8][1] , \data_i[8][0] , \data_i[7][31] ,
         \data_i[7][30] , \data_i[7][29] , \data_i[7][28] , \data_i[7][27] ,
         \data_i[7][26] , \data_i[7][25] , \data_i[7][24] , \data_i[7][23] ,
         \data_i[7][22] , \data_i[7][21] , \data_i[7][20] , \data_i[7][19] ,
         \data_i[7][18] , \data_i[7][17] , \data_i[7][16] , \data_i[7][15] ,
         \data_i[7][14] , \data_i[7][13] , \data_i[7][12] , \data_i[7][11] ,
         \data_i[7][10] , \data_i[7][9] , \data_i[7][8] , \data_i[7][7] ,
         \data_i[7][6] , \data_i[7][5] , \data_i[7][4] , \data_i[7][3] ,
         \data_i[7][2] , \data_i[7][1] , \data_i[7][0] , \data_i[6][31] ,
         \data_i[6][30] , \data_i[6][29] , \data_i[6][28] , \data_i[6][27] ,
         \data_i[6][26] , \data_i[6][25] , \data_i[6][24] , \data_i[6][23] ,
         \data_i[6][22] , \data_i[6][21] , \data_i[6][20] , \data_i[6][19] ,
         \data_i[6][18] , \data_i[6][17] , \data_i[6][16] , \data_i[6][15] ,
         \data_i[6][14] , \data_i[6][13] , \data_i[6][12] , \data_i[6][11] ,
         \data_i[6][10] , \data_i[6][9] , \data_i[6][8] , \data_i[6][7] ,
         \data_i[6][6] , \data_i[6][5] , \data_i[6][4] , \data_i[6][3] ,
         \data_i[6][2] , \data_i[6][1] , \data_i[6][0] , \data_i[5][31] ,
         \data_i[5][30] , \data_i[5][29] , \data_i[5][28] , \data_i[5][27] ,
         \data_i[5][26] , \data_i[5][25] , \data_i[5][24] , \data_i[5][23] ,
         \data_i[5][22] , \data_i[5][21] , \data_i[5][20] , \data_i[5][19] ,
         \data_i[5][18] , \data_i[5][17] , \data_i[5][16] , \data_i[5][15] ,
         \data_i[5][14] , \data_i[5][13] , \data_i[5][12] , \data_i[5][11] ,
         \data_i[5][10] , \data_i[5][9] , \data_i[5][8] , \data_i[5][7] ,
         \data_i[5][6] , \data_i[5][5] , \data_i[5][4] , \data_i[5][3] ,
         \data_i[5][2] , \data_i[5][1] , \data_i[5][0] , \data_i[4][31] ,
         \data_i[4][30] , \data_i[4][29] , \data_i[4][28] , \data_i[4][27] ,
         \data_i[4][26] , \data_i[4][25] , \data_i[4][24] , \data_i[4][23] ,
         \data_i[4][22] , \data_i[4][21] , \data_i[4][20] , \data_i[4][19] ,
         \data_i[4][18] , \data_i[4][17] , \data_i[4][16] , \data_i[4][15] ,
         \data_i[4][14] , \data_i[4][13] , \data_i[4][12] , \data_i[4][11] ,
         \data_i[4][10] , \data_i[4][9] , \data_i[4][8] , \data_i[4][7] ,
         \data_i[4][6] , \data_i[4][5] , \data_i[4][4] , \data_i[4][3] ,
         \data_i[4][2] , \data_i[4][1] , \data_i[4][0] , \data_i[3][31] ,
         \data_i[3][30] , \data_i[3][29] , \data_i[3][28] , \data_i[3][27] ,
         \data_i[3][26] , \data_i[3][25] , \data_i[3][24] , \data_i[3][23] ,
         \data_i[3][22] , \data_i[3][21] , \data_i[3][20] , \data_i[3][19] ,
         \data_i[3][18] , \data_i[3][17] , \data_i[3][16] , \data_i[3][15] ,
         \data_i[3][14] , \data_i[3][13] , \data_i[3][12] , \data_i[3][11] ,
         \data_i[3][10] , \data_i[3][9] , \data_i[3][8] , \data_i[3][7] ,
         \data_i[3][6] , \data_i[3][5] , \data_i[3][4] , \data_i[3][3] ,
         \data_i[3][2] , \data_i[3][1] , \data_i[3][0] , \data_i[2][31] ,
         \data_i[2][30] , \data_i[2][29] , \data_i[2][28] , \data_i[2][27] ,
         \data_i[2][26] , \data_i[2][25] , \data_i[2][24] , \data_i[2][23] ,
         \data_i[2][22] , \data_i[2][21] , \data_i[2][20] , \data_i[2][19] ,
         \data_i[2][18] , \data_i[2][17] , \data_i[2][16] , \data_i[2][15] ,
         \data_i[2][14] , \data_i[2][13] , \data_i[2][12] , \data_i[2][11] ,
         \data_i[2][10] , \data_i[2][9] , \data_i[2][8] , \data_i[2][7] ,
         \data_i[2][6] , \data_i[2][5] , \data_i[2][4] , \data_i[2][3] ,
         \data_i[2][2] , \data_i[2][1] , \data_i[2][0] , \data_i[1][31] ,
         \data_i[1][30] , \data_i[1][29] , \data_i[1][28] , \data_i[1][27] ,
         \data_i[1][26] , \data_i[1][25] , \data_i[1][24] , \data_i[1][23] ,
         \data_i[1][22] , \data_i[1][21] , \data_i[1][20] , \data_i[1][19] ,
         \data_i[1][18] , \data_i[1][17] , \data_i[1][16] , \data_i[1][15] ,
         \data_i[1][14] , \data_i[1][13] , \data_i[1][12] , \data_i[1][11] ,
         \data_i[1][10] , \data_i[1][9] , \data_i[1][8] , \data_i[1][7] ,
         \data_i[1][6] , \data_i[1][5] , \data_i[1][4] , \data_i[1][3] ,
         \data_i[1][2] , \data_i[1][1] , \data_i[1][0] , \data_i[0][31] ,
         \data_i[0][30] , \data_i[0][29] , \data_i[0][28] , \data_i[0][27] ,
         \data_i[0][26] , \data_i[0][25] , \data_i[0][24] , \data_i[0][23] ,
         \data_i[0][22] , \data_i[0][21] , \data_i[0][20] , \data_i[0][19] ,
         \data_i[0][18] , \data_i[0][17] , \data_i[0][16] , \data_i[0][15] ,
         \data_i[0][14] , \data_i[0][13] , \data_i[0][12] , \data_i[0][11] ,
         \data_i[0][10] , \data_i[0][9] , \data_i[0][8] , \data_i[0][7] ,
         \data_i[0][6] , \data_i[0][5] , \data_i[0][4] , \data_i[0][3] ,
         \data_i[0][2] , \data_i[0][1] , \data_i[0][0] ;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128;

  GTECH_AND2 C9 ( .A(N32), .B(N33), .Z(N37) );
  GTECH_AND2 C10 ( .A(N34), .B(N35), .Z(N38) );
  GTECH_AND2 C11 ( .A(N37), .B(N38), .Z(N39) );
  GTECH_AND2 C12 ( .A(N39), .B(N36), .Z(N40) );
  GTECH_OR2 C14 ( .A(select_i[4]), .B(select_i[3]), .Z(N41) );
  GTECH_OR2 C15 ( .A(select_i[2]), .B(select_i[1]), .Z(N42) );
  GTECH_OR2 C16 ( .A(N41), .B(N42), .Z(N43) );
  GTECH_OR2 C17 ( .A(N43), .B(N36), .Z(N44) );
  GTECH_OR2 C21 ( .A(select_i[2]), .B(N35), .Z(N46) );
  GTECH_OR2 C22 ( .A(N41), .B(N46), .Z(N47) );
  GTECH_OR2 C23 ( .A(N47), .B(select_i[0]), .Z(N48) );
  GTECH_OR2 C30 ( .A(N47), .B(N36), .Z(N50) );
  GTECH_OR2 C34 ( .A(N34), .B(select_i[1]), .Z(N52) );
  GTECH_OR2 C35 ( .A(N41), .B(N52), .Z(N53) );
  GTECH_OR2 C36 ( .A(N53), .B(select_i[0]), .Z(N54) );
  GTECH_OR2 C43 ( .A(N53), .B(N36), .Z(N56) );
  GTECH_OR2 C48 ( .A(N34), .B(N35), .Z(N58) );
  GTECH_OR2 C49 ( .A(N41), .B(N58), .Z(N59) );
  GTECH_OR2 C50 ( .A(N59), .B(select_i[0]), .Z(N60) );
  GTECH_OR2 C58 ( .A(N59), .B(N36), .Z(N62) );
  GTECH_OR2 C61 ( .A(select_i[4]), .B(N33), .Z(N64) );
  GTECH_OR2 C63 ( .A(N64), .B(N42), .Z(N65) );
  GTECH_OR2 C64 ( .A(N65), .B(select_i[0]), .Z(N66) );
  GTECH_OR2 C71 ( .A(N65), .B(N36), .Z(N68) );
  GTECH_OR2 C77 ( .A(N64), .B(N46), .Z(N70) );
  GTECH_OR2 C78 ( .A(N70), .B(select_i[0]), .Z(N71) );
  GTECH_OR2 C86 ( .A(N70), .B(N36), .Z(N73) );
  GTECH_OR2 C92 ( .A(N64), .B(N52), .Z(N75) );
  GTECH_OR2 C93 ( .A(N75), .B(select_i[0]), .Z(N76) );
  GTECH_OR2 C101 ( .A(N75), .B(N36), .Z(N78) );
  GTECH_OR2 C108 ( .A(N64), .B(N58), .Z(N80) );
  GTECH_OR2 C109 ( .A(N80), .B(select_i[0]), .Z(N81) );
  GTECH_OR2 C118 ( .A(N80), .B(N36), .Z(N83) );
  GTECH_OR2 C121 ( .A(N32), .B(select_i[3]), .Z(N85) );
  GTECH_OR2 C123 ( .A(N85), .B(N42), .Z(N86) );
  GTECH_OR2 C124 ( .A(N86), .B(select_i[0]), .Z(N87) );
  GTECH_OR2 C131 ( .A(N86), .B(N36), .Z(N89) );
  GTECH_OR2 C137 ( .A(N85), .B(N46), .Z(N91) );
  GTECH_OR2 C138 ( .A(N91), .B(select_i[0]), .Z(N92) );
  GTECH_OR2 C146 ( .A(N91), .B(N36), .Z(N94) );
  GTECH_OR2 C152 ( .A(N85), .B(N52), .Z(N96) );
  GTECH_OR2 C153 ( .A(N96), .B(select_i[0]), .Z(N97) );
  GTECH_OR2 C161 ( .A(N96), .B(N36), .Z(N99) );
  GTECH_OR2 C168 ( .A(N85), .B(N58), .Z(N101) );
  GTECH_OR2 C169 ( .A(N101), .B(select_i[0]), .Z(N102) );
  GTECH_OR2 C178 ( .A(N101), .B(N36), .Z(N104) );
  GTECH_OR2 C182 ( .A(N32), .B(N33), .Z(N106) );
  GTECH_OR2 C184 ( .A(N106), .B(N42), .Z(N107) );
  GTECH_OR2 C185 ( .A(N107), .B(select_i[0]), .Z(N108) );
  GTECH_OR2 C193 ( .A(N107), .B(N36), .Z(N110) );
  GTECH_OR2 C200 ( .A(N106), .B(N46), .Z(N112) );
  GTECH_OR2 C201 ( .A(N112), .B(select_i[0]), .Z(N113) );
  GTECH_OR2 C210 ( .A(N112), .B(N36), .Z(N115) );
  GTECH_OR2 C217 ( .A(N106), .B(N52), .Z(N117) );
  GTECH_OR2 C218 ( .A(N117), .B(select_i[0]), .Z(N118) );
  GTECH_OR2 C227 ( .A(N117), .B(N36), .Z(N120) );
  GTECH_OR2 C235 ( .A(N106), .B(N58), .Z(N122) );
  GTECH_OR2 C236 ( .A(N122), .B(select_i[0]), .Z(N123) );
  GTECH_AND2 C238 ( .A(select_i[4]), .B(select_i[3]), .Z(N125) );
  GTECH_AND2 C239 ( .A(select_i[2]), .B(select_i[1]), .Z(N126) );
  GTECH_AND2 C240 ( .A(N125), .B(N126), .Z(N127) );
  GTECH_AND2 C241 ( .A(N127), .B(select_i[0]), .Z(N128) );
  SELECT_OP C339 ( .DATA1({\data_i[0][31] , \data_i[0][30] , \data_i[0][29] , 
        \data_i[0][28] , \data_i[0][27] , \data_i[0][26] , \data_i[0][25] , 
        \data_i[0][24] , \data_i[0][23] , \data_i[0][22] , \data_i[0][21] , 
        \data_i[0][20] , \data_i[0][19] , \data_i[0][18] , \data_i[0][17] , 
        \data_i[0][16] , \data_i[0][15] , \data_i[0][14] , \data_i[0][13] , 
        \data_i[0][12] , \data_i[0][11] , \data_i[0][10] , \data_i[0][9] , 
        \data_i[0][8] , \data_i[0][7] , \data_i[0][6] , \data_i[0][5] , 
        \data_i[0][4] , \data_i[0][3] , \data_i[0][2] , \data_i[0][1] , 
        \data_i[0][0] }), .DATA2({\data_i[1][31] , \data_i[1][30] , 
        \data_i[1][29] , \data_i[1][28] , \data_i[1][27] , \data_i[1][26] , 
        \data_i[1][25] , \data_i[1][24] , \data_i[1][23] , \data_i[1][22] , 
        \data_i[1][21] , \data_i[1][20] , \data_i[1][19] , \data_i[1][18] , 
        \data_i[1][17] , \data_i[1][16] , \data_i[1][15] , \data_i[1][14] , 
        \data_i[1][13] , \data_i[1][12] , \data_i[1][11] , \data_i[1][10] , 
        \data_i[1][9] , \data_i[1][8] , \data_i[1][7] , \data_i[1][6] , 
        \data_i[1][5] , \data_i[1][4] , \data_i[1][3] , \data_i[1][2] , 
        \data_i[1][1] , \data_i[1][0] }), .DATA3({\data_i[2][31] , 
        \data_i[2][30] , \data_i[2][29] , \data_i[2][28] , \data_i[2][27] , 
        \data_i[2][26] , \data_i[2][25] , \data_i[2][24] , \data_i[2][23] , 
        \data_i[2][22] , \data_i[2][21] , \data_i[2][20] , \data_i[2][19] , 
        \data_i[2][18] , \data_i[2][17] , \data_i[2][16] , \data_i[2][15] , 
        \data_i[2][14] , \data_i[2][13] , \data_i[2][12] , \data_i[2][11] , 
        \data_i[2][10] , \data_i[2][9] , \data_i[2][8] , \data_i[2][7] , 
        \data_i[2][6] , \data_i[2][5] , \data_i[2][4] , \data_i[2][3] , 
        \data_i[2][2] , \data_i[2][1] , \data_i[2][0] }), .DATA4({
        \data_i[3][31] , \data_i[3][30] , \data_i[3][29] , \data_i[3][28] , 
        \data_i[3][27] , \data_i[3][26] , \data_i[3][25] , \data_i[3][24] , 
        \data_i[3][23] , \data_i[3][22] , \data_i[3][21] , \data_i[3][20] , 
        \data_i[3][19] , \data_i[3][18] , \data_i[3][17] , \data_i[3][16] , 
        \data_i[3][15] , \data_i[3][14] , \data_i[3][13] , \data_i[3][12] , 
        \data_i[3][11] , \data_i[3][10] , \data_i[3][9] , \data_i[3][8] , 
        \data_i[3][7] , \data_i[3][6] , \data_i[3][5] , \data_i[3][4] , 
        \data_i[3][3] , \data_i[3][2] , \data_i[3][1] , \data_i[3][0] }), 
        .DATA5({\data_i[4][31] , \data_i[4][30] , \data_i[4][29] , 
        \data_i[4][28] , \data_i[4][27] , \data_i[4][26] , \data_i[4][25] , 
        \data_i[4][24] , \data_i[4][23] , \data_i[4][22] , \data_i[4][21] , 
        \data_i[4][20] , \data_i[4][19] , \data_i[4][18] , \data_i[4][17] , 
        \data_i[4][16] , \data_i[4][15] , \data_i[4][14] , \data_i[4][13] , 
        \data_i[4][12] , \data_i[4][11] , \data_i[4][10] , \data_i[4][9] , 
        \data_i[4][8] , \data_i[4][7] , \data_i[4][6] , \data_i[4][5] , 
        \data_i[4][4] , \data_i[4][3] , \data_i[4][2] , \data_i[4][1] , 
        \data_i[4][0] }), .DATA6({\data_i[5][31] , \data_i[5][30] , 
        \data_i[5][29] , \data_i[5][28] , \data_i[5][27] , \data_i[5][26] , 
        \data_i[5][25] , \data_i[5][24] , \data_i[5][23] , \data_i[5][22] , 
        \data_i[5][21] , \data_i[5][20] , \data_i[5][19] , \data_i[5][18] , 
        \data_i[5][17] , \data_i[5][16] , \data_i[5][15] , \data_i[5][14] , 
        \data_i[5][13] , \data_i[5][12] , \data_i[5][11] , \data_i[5][10] , 
        \data_i[5][9] , \data_i[5][8] , \data_i[5][7] , \data_i[5][6] , 
        \data_i[5][5] , \data_i[5][4] , \data_i[5][3] , \data_i[5][2] , 
        \data_i[5][1] , \data_i[5][0] }), .DATA7({\data_i[6][31] , 
        \data_i[6][30] , \data_i[6][29] , \data_i[6][28] , \data_i[6][27] , 
        \data_i[6][26] , \data_i[6][25] , \data_i[6][24] , \data_i[6][23] , 
        \data_i[6][22] , \data_i[6][21] , \data_i[6][20] , \data_i[6][19] , 
        \data_i[6][18] , \data_i[6][17] , \data_i[6][16] , \data_i[6][15] , 
        \data_i[6][14] , \data_i[6][13] , \data_i[6][12] , \data_i[6][11] , 
        \data_i[6][10] , \data_i[6][9] , \data_i[6][8] , \data_i[6][7] , 
        \data_i[6][6] , \data_i[6][5] , \data_i[6][4] , \data_i[6][3] , 
        \data_i[6][2] , \data_i[6][1] , \data_i[6][0] }), .DATA8({
        \data_i[7][31] , \data_i[7][30] , \data_i[7][29] , \data_i[7][28] , 
        \data_i[7][27] , \data_i[7][26] , \data_i[7][25] , \data_i[7][24] , 
        \data_i[7][23] , \data_i[7][22] , \data_i[7][21] , \data_i[7][20] , 
        \data_i[7][19] , \data_i[7][18] , \data_i[7][17] , \data_i[7][16] , 
        \data_i[7][15] , \data_i[7][14] , \data_i[7][13] , \data_i[7][12] , 
        \data_i[7][11] , \data_i[7][10] , \data_i[7][9] , \data_i[7][8] , 
        \data_i[7][7] , \data_i[7][6] , \data_i[7][5] , \data_i[7][4] , 
        \data_i[7][3] , \data_i[7][2] , \data_i[7][1] , \data_i[7][0] }), 
        .DATA9({\data_i[8][31] , \data_i[8][30] , \data_i[8][29] , 
        \data_i[8][28] , \data_i[8][27] , \data_i[8][26] , \data_i[8][25] , 
        \data_i[8][24] , \data_i[8][23] , \data_i[8][22] , \data_i[8][21] , 
        \data_i[8][20] , \data_i[8][19] , \data_i[8][18] , \data_i[8][17] , 
        \data_i[8][16] , \data_i[8][15] , \data_i[8][14] , \data_i[8][13] , 
        \data_i[8][12] , \data_i[8][11] , \data_i[8][10] , \data_i[8][9] , 
        \data_i[8][8] , \data_i[8][7] , \data_i[8][6] , \data_i[8][5] , 
        \data_i[8][4] , \data_i[8][3] , \data_i[8][2] , \data_i[8][1] , 
        \data_i[8][0] }), .DATA10({\data_i[9][31] , \data_i[9][30] , 
        \data_i[9][29] , \data_i[9][28] , \data_i[9][27] , \data_i[9][26] , 
        \data_i[9][25] , \data_i[9][24] , \data_i[9][23] , \data_i[9][22] , 
        \data_i[9][21] , \data_i[9][20] , \data_i[9][19] , \data_i[9][18] , 
        \data_i[9][17] , \data_i[9][16] , \data_i[9][15] , \data_i[9][14] , 
        \data_i[9][13] , \data_i[9][12] , \data_i[9][11] , \data_i[9][10] , 
        \data_i[9][9] , \data_i[9][8] , \data_i[9][7] , \data_i[9][6] , 
        \data_i[9][5] , \data_i[9][4] , \data_i[9][3] , \data_i[9][2] , 
        \data_i[9][1] , \data_i[9][0] }), .DATA11({\data_i[10][31] , 
        \data_i[10][30] , \data_i[10][29] , \data_i[10][28] , \data_i[10][27] , 
        \data_i[10][26] , \data_i[10][25] , \data_i[10][24] , \data_i[10][23] , 
        \data_i[10][22] , \data_i[10][21] , \data_i[10][20] , \data_i[10][19] , 
        \data_i[10][18] , \data_i[10][17] , \data_i[10][16] , \data_i[10][15] , 
        \data_i[10][14] , \data_i[10][13] , \data_i[10][12] , \data_i[10][11] , 
        \data_i[10][10] , \data_i[10][9] , \data_i[10][8] , \data_i[10][7] , 
        \data_i[10][6] , \data_i[10][5] , \data_i[10][4] , \data_i[10][3] , 
        \data_i[10][2] , \data_i[10][1] , \data_i[10][0] }), .DATA12({
        \data_i[11][31] , \data_i[11][30] , \data_i[11][29] , \data_i[11][28] , 
        \data_i[11][27] , \data_i[11][26] , \data_i[11][25] , \data_i[11][24] , 
        \data_i[11][23] , \data_i[11][22] , \data_i[11][21] , \data_i[11][20] , 
        \data_i[11][19] , \data_i[11][18] , \data_i[11][17] , \data_i[11][16] , 
        \data_i[11][15] , \data_i[11][14] , \data_i[11][13] , \data_i[11][12] , 
        \data_i[11][11] , \data_i[11][10] , \data_i[11][9] , \data_i[11][8] , 
        \data_i[11][7] , \data_i[11][6] , \data_i[11][5] , \data_i[11][4] , 
        \data_i[11][3] , \data_i[11][2] , \data_i[11][1] , \data_i[11][0] }), 
        .DATA13({\data_i[12][31] , \data_i[12][30] , \data_i[12][29] , 
        \data_i[12][28] , \data_i[12][27] , \data_i[12][26] , \data_i[12][25] , 
        \data_i[12][24] , \data_i[12][23] , \data_i[12][22] , \data_i[12][21] , 
        \data_i[12][20] , \data_i[12][19] , \data_i[12][18] , \data_i[12][17] , 
        \data_i[12][16] , \data_i[12][15] , \data_i[12][14] , \data_i[12][13] , 
        \data_i[12][12] , \data_i[12][11] , \data_i[12][10] , \data_i[12][9] , 
        \data_i[12][8] , \data_i[12][7] , \data_i[12][6] , \data_i[12][5] , 
        \data_i[12][4] , \data_i[12][3] , \data_i[12][2] , \data_i[12][1] , 
        \data_i[12][0] }), .DATA14({\data_i[13][31] , \data_i[13][30] , 
        \data_i[13][29] , \data_i[13][28] , \data_i[13][27] , \data_i[13][26] , 
        \data_i[13][25] , \data_i[13][24] , \data_i[13][23] , \data_i[13][22] , 
        \data_i[13][21] , \data_i[13][20] , \data_i[13][19] , \data_i[13][18] , 
        \data_i[13][17] , \data_i[13][16] , \data_i[13][15] , \data_i[13][14] , 
        \data_i[13][13] , \data_i[13][12] , \data_i[13][11] , \data_i[13][10] , 
        \data_i[13][9] , \data_i[13][8] , \data_i[13][7] , \data_i[13][6] , 
        \data_i[13][5] , \data_i[13][4] , \data_i[13][3] , \data_i[13][2] , 
        \data_i[13][1] , \data_i[13][0] }), .DATA15({\data_i[14][31] , 
        \data_i[14][30] , \data_i[14][29] , \data_i[14][28] , \data_i[14][27] , 
        \data_i[14][26] , \data_i[14][25] , \data_i[14][24] , \data_i[14][23] , 
        \data_i[14][22] , \data_i[14][21] , \data_i[14][20] , \data_i[14][19] , 
        \data_i[14][18] , \data_i[14][17] , \data_i[14][16] , \data_i[14][15] , 
        \data_i[14][14] , \data_i[14][13] , \data_i[14][12] , \data_i[14][11] , 
        \data_i[14][10] , \data_i[14][9] , \data_i[14][8] , \data_i[14][7] , 
        \data_i[14][6] , \data_i[14][5] , \data_i[14][4] , \data_i[14][3] , 
        \data_i[14][2] , \data_i[14][1] , \data_i[14][0] }), .DATA16({
        \data_i[15][31] , \data_i[15][30] , \data_i[15][29] , \data_i[15][28] , 
        \data_i[15][27] , \data_i[15][26] , \data_i[15][25] , \data_i[15][24] , 
        \data_i[15][23] , \data_i[15][22] , \data_i[15][21] , \data_i[15][20] , 
        \data_i[15][19] , \data_i[15][18] , \data_i[15][17] , \data_i[15][16] , 
        \data_i[15][15] , \data_i[15][14] , \data_i[15][13] , \data_i[15][12] , 
        \data_i[15][11] , \data_i[15][10] , \data_i[15][9] , \data_i[15][8] , 
        \data_i[15][7] , \data_i[15][6] , \data_i[15][5] , \data_i[15][4] , 
        \data_i[15][3] , \data_i[15][2] , \data_i[15][1] , \data_i[15][0] }), 
        .DATA17({\data_i[16][31] , \data_i[16][30] , \data_i[16][29] , 
        \data_i[16][28] , \data_i[16][27] , \data_i[16][26] , \data_i[16][25] , 
        \data_i[16][24] , \data_i[16][23] , \data_i[16][22] , \data_i[16][21] , 
        \data_i[16][20] , \data_i[16][19] , \data_i[16][18] , \data_i[16][17] , 
        \data_i[16][16] , \data_i[16][15] , \data_i[16][14] , \data_i[16][13] , 
        \data_i[16][12] , \data_i[16][11] , \data_i[16][10] , \data_i[16][9] , 
        \data_i[16][8] , \data_i[16][7] , \data_i[16][6] , \data_i[16][5] , 
        \data_i[16][4] , \data_i[16][3] , \data_i[16][2] , \data_i[16][1] , 
        \data_i[16][0] }), .DATA18({\data_i[17][31] , \data_i[17][30] , 
        \data_i[17][29] , \data_i[17][28] , \data_i[17][27] , \data_i[17][26] , 
        \data_i[17][25] , \data_i[17][24] , \data_i[17][23] , \data_i[17][22] , 
        \data_i[17][21] , \data_i[17][20] , \data_i[17][19] , \data_i[17][18] , 
        \data_i[17][17] , \data_i[17][16] , \data_i[17][15] , \data_i[17][14] , 
        \data_i[17][13] , \data_i[17][12] , \data_i[17][11] , \data_i[17][10] , 
        \data_i[17][9] , \data_i[17][8] , \data_i[17][7] , \data_i[17][6] , 
        \data_i[17][5] , \data_i[17][4] , \data_i[17][3] , \data_i[17][2] , 
        \data_i[17][1] , \data_i[17][0] }), .DATA19({\data_i[18][31] , 
        \data_i[18][30] , \data_i[18][29] , \data_i[18][28] , \data_i[18][27] , 
        \data_i[18][26] , \data_i[18][25] , \data_i[18][24] , \data_i[18][23] , 
        \data_i[18][22] , \data_i[18][21] , \data_i[18][20] , \data_i[18][19] , 
        \data_i[18][18] , \data_i[18][17] , \data_i[18][16] , \data_i[18][15] , 
        \data_i[18][14] , \data_i[18][13] , \data_i[18][12] , \data_i[18][11] , 
        \data_i[18][10] , \data_i[18][9] , \data_i[18][8] , \data_i[18][7] , 
        \data_i[18][6] , \data_i[18][5] , \data_i[18][4] , \data_i[18][3] , 
        \data_i[18][2] , \data_i[18][1] , \data_i[18][0] }), .DATA20({
        \data_i[19][31] , \data_i[19][30] , \data_i[19][29] , \data_i[19][28] , 
        \data_i[19][27] , \data_i[19][26] , \data_i[19][25] , \data_i[19][24] , 
        \data_i[19][23] , \data_i[19][22] , \data_i[19][21] , \data_i[19][20] , 
        \data_i[19][19] , \data_i[19][18] , \data_i[19][17] , \data_i[19][16] , 
        \data_i[19][15] , \data_i[19][14] , \data_i[19][13] , \data_i[19][12] , 
        \data_i[19][11] , \data_i[19][10] , \data_i[19][9] , \data_i[19][8] , 
        \data_i[19][7] , \data_i[19][6] , \data_i[19][5] , \data_i[19][4] , 
        \data_i[19][3] , \data_i[19][2] , \data_i[19][1] , \data_i[19][0] }), 
        .DATA21({\data_i[20][31] , \data_i[20][30] , \data_i[20][29] , 
        \data_i[20][28] , \data_i[20][27] , \data_i[20][26] , \data_i[20][25] , 
        \data_i[20][24] , \data_i[20][23] , \data_i[20][22] , \data_i[20][21] , 
        \data_i[20][20] , \data_i[20][19] , \data_i[20][18] , \data_i[20][17] , 
        \data_i[20][16] , \data_i[20][15] , \data_i[20][14] , \data_i[20][13] , 
        \data_i[20][12] , \data_i[20][11] , \data_i[20][10] , \data_i[20][9] , 
        \data_i[20][8] , \data_i[20][7] , \data_i[20][6] , \data_i[20][5] , 
        \data_i[20][4] , \data_i[20][3] , \data_i[20][2] , \data_i[20][1] , 
        \data_i[20][0] }), .DATA22({\data_i[21][31] , \data_i[21][30] , 
        \data_i[21][29] , \data_i[21][28] , \data_i[21][27] , \data_i[21][26] , 
        \data_i[21][25] , \data_i[21][24] , \data_i[21][23] , \data_i[21][22] , 
        \data_i[21][21] , \data_i[21][20] , \data_i[21][19] , \data_i[21][18] , 
        \data_i[21][17] , \data_i[21][16] , \data_i[21][15] , \data_i[21][14] , 
        \data_i[21][13] , \data_i[21][12] , \data_i[21][11] , \data_i[21][10] , 
        \data_i[21][9] , \data_i[21][8] , \data_i[21][7] , \data_i[21][6] , 
        \data_i[21][5] , \data_i[21][4] , \data_i[21][3] , \data_i[21][2] , 
        \data_i[21][1] , \data_i[21][0] }), .DATA23({\data_i[22][31] , 
        \data_i[22][30] , \data_i[22][29] , \data_i[22][28] , \data_i[22][27] , 
        \data_i[22][26] , \data_i[22][25] , \data_i[22][24] , \data_i[22][23] , 
        \data_i[22][22] , \data_i[22][21] , \data_i[22][20] , \data_i[22][19] , 
        \data_i[22][18] , \data_i[22][17] , \data_i[22][16] , \data_i[22][15] , 
        \data_i[22][14] , \data_i[22][13] , \data_i[22][12] , \data_i[22][11] , 
        \data_i[22][10] , \data_i[22][9] , \data_i[22][8] , \data_i[22][7] , 
        \data_i[22][6] , \data_i[22][5] , \data_i[22][4] , \data_i[22][3] , 
        \data_i[22][2] , \data_i[22][1] , \data_i[22][0] }), .DATA24({
        \data_i[23][31] , \data_i[23][30] , \data_i[23][29] , \data_i[23][28] , 
        \data_i[23][27] , \data_i[23][26] , \data_i[23][25] , \data_i[23][24] , 
        \data_i[23][23] , \data_i[23][22] , \data_i[23][21] , \data_i[23][20] , 
        \data_i[23][19] , \data_i[23][18] , \data_i[23][17] , \data_i[23][16] , 
        \data_i[23][15] , \data_i[23][14] , \data_i[23][13] , \data_i[23][12] , 
        \data_i[23][11] , \data_i[23][10] , \data_i[23][9] , \data_i[23][8] , 
        \data_i[23][7] , \data_i[23][6] , \data_i[23][5] , \data_i[23][4] , 
        \data_i[23][3] , \data_i[23][2] , \data_i[23][1] , \data_i[23][0] }), 
        .DATA25({\data_i[24][31] , \data_i[24][30] , \data_i[24][29] , 
        \data_i[24][28] , \data_i[24][27] , \data_i[24][26] , \data_i[24][25] , 
        \data_i[24][24] , \data_i[24][23] , \data_i[24][22] , \data_i[24][21] , 
        \data_i[24][20] , \data_i[24][19] , \data_i[24][18] , \data_i[24][17] , 
        \data_i[24][16] , \data_i[24][15] , \data_i[24][14] , \data_i[24][13] , 
        \data_i[24][12] , \data_i[24][11] , \data_i[24][10] , \data_i[24][9] , 
        \data_i[24][8] , \data_i[24][7] , \data_i[24][6] , \data_i[24][5] , 
        \data_i[24][4] , \data_i[24][3] , \data_i[24][2] , \data_i[24][1] , 
        \data_i[24][0] }), .DATA26({\data_i[25][31] , \data_i[25][30] , 
        \data_i[25][29] , \data_i[25][28] , \data_i[25][27] , \data_i[25][26] , 
        \data_i[25][25] , \data_i[25][24] , \data_i[25][23] , \data_i[25][22] , 
        \data_i[25][21] , \data_i[25][20] , \data_i[25][19] , \data_i[25][18] , 
        \data_i[25][17] , \data_i[25][16] , \data_i[25][15] , \data_i[25][14] , 
        \data_i[25][13] , \data_i[25][12] , \data_i[25][11] , \data_i[25][10] , 
        \data_i[25][9] , \data_i[25][8] , \data_i[25][7] , \data_i[25][6] , 
        \data_i[25][5] , \data_i[25][4] , \data_i[25][3] , \data_i[25][2] , 
        \data_i[25][1] , \data_i[25][0] }), .DATA27({\data_i[26][31] , 
        \data_i[26][30] , \data_i[26][29] , \data_i[26][28] , \data_i[26][27] , 
        \data_i[26][26] , \data_i[26][25] , \data_i[26][24] , \data_i[26][23] , 
        \data_i[26][22] , \data_i[26][21] , \data_i[26][20] , \data_i[26][19] , 
        \data_i[26][18] , \data_i[26][17] , \data_i[26][16] , \data_i[26][15] , 
        \data_i[26][14] , \data_i[26][13] , \data_i[26][12] , \data_i[26][11] , 
        \data_i[26][10] , \data_i[26][9] , \data_i[26][8] , \data_i[26][7] , 
        \data_i[26][6] , \data_i[26][5] , \data_i[26][4] , \data_i[26][3] , 
        \data_i[26][2] , \data_i[26][1] , \data_i[26][0] }), .DATA28({
        \data_i[27][31] , \data_i[27][30] , \data_i[27][29] , \data_i[27][28] , 
        \data_i[27][27] , \data_i[27][26] , \data_i[27][25] , \data_i[27][24] , 
        \data_i[27][23] , \data_i[27][22] , \data_i[27][21] , \data_i[27][20] , 
        \data_i[27][19] , \data_i[27][18] , \data_i[27][17] , \data_i[27][16] , 
        \data_i[27][15] , \data_i[27][14] , \data_i[27][13] , \data_i[27][12] , 
        \data_i[27][11] , \data_i[27][10] , \data_i[27][9] , \data_i[27][8] , 
        \data_i[27][7] , \data_i[27][6] , \data_i[27][5] , \data_i[27][4] , 
        \data_i[27][3] , \data_i[27][2] , \data_i[27][1] , \data_i[27][0] }), 
        .DATA29({\data_i[28][31] , \data_i[28][30] , \data_i[28][29] , 
        \data_i[28][28] , \data_i[28][27] , \data_i[28][26] , \data_i[28][25] , 
        \data_i[28][24] , \data_i[28][23] , \data_i[28][22] , \data_i[28][21] , 
        \data_i[28][20] , \data_i[28][19] , \data_i[28][18] , \data_i[28][17] , 
        \data_i[28][16] , \data_i[28][15] , \data_i[28][14] , \data_i[28][13] , 
        \data_i[28][12] , \data_i[28][11] , \data_i[28][10] , \data_i[28][9] , 
        \data_i[28][8] , \data_i[28][7] , \data_i[28][6] , \data_i[28][5] , 
        \data_i[28][4] , \data_i[28][3] , \data_i[28][2] , \data_i[28][1] , 
        \data_i[28][0] }), .DATA30({\data_i[29][31] , \data_i[29][30] , 
        \data_i[29][29] , \data_i[29][28] , \data_i[29][27] , \data_i[29][26] , 
        \data_i[29][25] , \data_i[29][24] , \data_i[29][23] , \data_i[29][22] , 
        \data_i[29][21] , \data_i[29][20] , \data_i[29][19] , \data_i[29][18] , 
        \data_i[29][17] , \data_i[29][16] , \data_i[29][15] , \data_i[29][14] , 
        \data_i[29][13] , \data_i[29][12] , \data_i[29][11] , \data_i[29][10] , 
        \data_i[29][9] , \data_i[29][8] , \data_i[29][7] , \data_i[29][6] , 
        \data_i[29][5] , \data_i[29][4] , \data_i[29][3] , \data_i[29][2] , 
        \data_i[29][1] , \data_i[29][0] }), .DATA31({\data_i[30][31] , 
        \data_i[30][30] , \data_i[30][29] , \data_i[30][28] , \data_i[30][27] , 
        \data_i[30][26] , \data_i[30][25] , \data_i[30][24] , \data_i[30][23] , 
        \data_i[30][22] , \data_i[30][21] , \data_i[30][20] , \data_i[30][19] , 
        \data_i[30][18] , \data_i[30][17] , \data_i[30][16] , \data_i[30][15] , 
        \data_i[30][14] , \data_i[30][13] , \data_i[30][12] , \data_i[30][11] , 
        \data_i[30][10] , \data_i[30][9] , \data_i[30][8] , \data_i[30][7] , 
        \data_i[30][6] , \data_i[30][5] , \data_i[30][4] , \data_i[30][3] , 
        \data_i[30][2] , \data_i[30][1] , \data_i[30][0] }), .DATA32({
        \data_i[31][31] , \data_i[31][30] , \data_i[31][29] , \data_i[31][28] , 
        \data_i[31][27] , \data_i[31][26] , \data_i[31][25] , \data_i[31][24] , 
        \data_i[31][23] , \data_i[31][22] , \data_i[31][21] , \data_i[31][20] , 
        \data_i[31][19] , \data_i[31][18] , \data_i[31][17] , \data_i[31][16] , 
        \data_i[31][15] , \data_i[31][14] , \data_i[31][13] , \data_i[31][12] , 
        \data_i[31][11] , \data_i[31][10] , \data_i[31][9] , \data_i[31][8] , 
        \data_i[31][7] , \data_i[31][6] , \data_i[31][5] , \data_i[31][4] , 
        \data_i[31][3] , \data_i[31][2] , \data_i[31][1] , \data_i[31][0] }), 
        .CONTROL1(N0), .CONTROL2(N1), .CONTROL3(N2), .CONTROL4(N3), .CONTROL5(
        N4), .CONTROL6(N5), .CONTROL7(N6), .CONTROL8(N7), .CONTROL9(N8), 
        .CONTROL10(N9), .CONTROL11(N10), .CONTROL12(N11), .CONTROL13(N12), 
        .CONTROL14(N13), .CONTROL15(N14), .CONTROL16(N15), .CONTROL17(N16), 
        .CONTROL18(N17), .CONTROL19(N18), .CONTROL20(N19), .CONTROL21(N20), 
        .CONTROL22(N21), .CONTROL23(N22), .CONTROL24(N23), .CONTROL25(N24), 
        .CONTROL26(N25), .CONTROL27(N26), .CONTROL28(N27), .CONTROL29(N28), 
        .CONTROL30(N29), .CONTROL31(N30), .CONTROL32(N31), .Z(data_o) );
  GTECH_BUF B_0 ( .A(N40), .Z(N0) );
  GTECH_BUF B_1 ( .A(N45), .Z(N1) );
  GTECH_BUF B_2 ( .A(N49), .Z(N2) );
  GTECH_BUF B_3 ( .A(N51), .Z(N3) );
  GTECH_BUF B_4 ( .A(N55), .Z(N4) );
  GTECH_BUF B_5 ( .A(N57), .Z(N5) );
  GTECH_BUF B_6 ( .A(N61), .Z(N6) );
  GTECH_BUF B_7 ( .A(N63), .Z(N7) );
  GTECH_BUF B_8 ( .A(N67), .Z(N8) );
  GTECH_BUF B_9 ( .A(N69), .Z(N9) );
  GTECH_BUF B_10 ( .A(N72), .Z(N10) );
  GTECH_BUF B_11 ( .A(N74), .Z(N11) );
  GTECH_BUF B_12 ( .A(N77), .Z(N12) );
  GTECH_BUF B_13 ( .A(N79), .Z(N13) );
  GTECH_BUF B_14 ( .A(N82), .Z(N14) );
  GTECH_BUF B_15 ( .A(N84), .Z(N15) );
  GTECH_BUF B_16 ( .A(N88), .Z(N16) );
  GTECH_BUF B_17 ( .A(N90), .Z(N17) );
  GTECH_BUF B_18 ( .A(N93), .Z(N18) );
  GTECH_BUF B_19 ( .A(N95), .Z(N19) );
  GTECH_BUF B_20 ( .A(N98), .Z(N20) );
  GTECH_BUF B_21 ( .A(N100), .Z(N21) );
  GTECH_BUF B_22 ( .A(N103), .Z(N22) );
  GTECH_BUF B_23 ( .A(N105), .Z(N23) );
  GTECH_BUF B_24 ( .A(N109), .Z(N24) );
  GTECH_BUF B_25 ( .A(N111), .Z(N25) );
  GTECH_BUF B_26 ( .A(N114), .Z(N26) );
  GTECH_BUF B_27 ( .A(N116), .Z(N27) );
  GTECH_BUF B_28 ( .A(N119), .Z(N28) );
  GTECH_BUF B_29 ( .A(N121), .Z(N29) );
  GTECH_BUF B_30 ( .A(N124), .Z(N30) );
  GTECH_BUF B_31 ( .A(N128), .Z(N31) );
  GTECH_NOT I_0 ( .A(select_i[4]), .Z(N32) );
  GTECH_NOT I_1 ( .A(select_i[3]), .Z(N33) );
  GTECH_NOT I_2 ( .A(select_i[2]), .Z(N34) );
  GTECH_NOT I_3 ( .A(select_i[1]), .Z(N35) );
  GTECH_NOT I_4 ( .A(select_i[0]), .Z(N36) );
  GTECH_NOT I_5 ( .A(N44), .Z(N45) );
  GTECH_NOT I_6 ( .A(N48), .Z(N49) );
  GTECH_NOT I_7 ( .A(N50), .Z(N51) );
  GTECH_NOT I_8 ( .A(N54), .Z(N55) );
  GTECH_NOT I_9 ( .A(N56), .Z(N57) );
  GTECH_NOT I_10 ( .A(N60), .Z(N61) );
  GTECH_NOT I_11 ( .A(N62), .Z(N63) );
  GTECH_NOT I_12 ( .A(N66), .Z(N67) );
  GTECH_NOT I_13 ( .A(N68), .Z(N69) );
  GTECH_NOT I_14 ( .A(N71), .Z(N72) );
  GTECH_NOT I_15 ( .A(N73), .Z(N74) );
  GTECH_NOT I_16 ( .A(N76), .Z(N77) );
  GTECH_NOT I_17 ( .A(N78), .Z(N79) );
  GTECH_NOT I_18 ( .A(N81), .Z(N82) );
  GTECH_NOT I_19 ( .A(N83), .Z(N84) );
  GTECH_NOT I_20 ( .A(N87), .Z(N88) );
  GTECH_NOT I_21 ( .A(N89), .Z(N90) );
  GTECH_NOT I_22 ( .A(N92), .Z(N93) );
  GTECH_NOT I_23 ( .A(N94), .Z(N95) );
  GTECH_NOT I_24 ( .A(N97), .Z(N98) );
  GTECH_NOT I_25 ( .A(N99), .Z(N100) );
  GTECH_NOT I_26 ( .A(N102), .Z(N103) );
  GTECH_NOT I_27 ( .A(N104), .Z(N105) );
  GTECH_NOT I_28 ( .A(N108), .Z(N109) );
  GTECH_NOT I_29 ( .A(N110), .Z(N111) );
  GTECH_NOT I_30 ( .A(N113), .Z(N114) );
  GTECH_NOT I_31 ( .A(N115), .Z(N116) );
  GTECH_NOT I_32 ( .A(N118), .Z(N119) );
  GTECH_NOT I_33 ( .A(N120), .Z(N121) );
  GTECH_NOT I_34 ( .A(N123), .Z(N124) );
endmodule


module FF_WIDTH32_31 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_31 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_31 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_31 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_31 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_0 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_0 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_0 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_0 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_0 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_1 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_1 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_1 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_1 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_1 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_2 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_2 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_2 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_2 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_2 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_3 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_3 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_3 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_3 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_3 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_4 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_4 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_4 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_4 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_4 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_5 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_5 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_5 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_5 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_5 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_6 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_6 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_6 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_6 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_6 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_7 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_7 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_7 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_7 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_7 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_8 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_8 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_8 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_8 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_8 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_9 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_9 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_9 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_9 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_9 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_10 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_10 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_10 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_10 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_10 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_11 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_11 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_11 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_11 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_11 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_12 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_12 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_12 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_12 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_12 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_13 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_13 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_13 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_13 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_13 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_14 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_14 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_14 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_14 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_14 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_15 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_15 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_15 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_15 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_15 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_16 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_16 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_16 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_16 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_16 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_17 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_17 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_17 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_17 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_17 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_18 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_18 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_18 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_18 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_18 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_19 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_19 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_19 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_19 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_19 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_20 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_20 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_20 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_20 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_20 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_21 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_21 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_21 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_21 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_21 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_22 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_22 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_22 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_22 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_22 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_23 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_23 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_23 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_23 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_23 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_24 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_24 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_24 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_24 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_24 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_25 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_25 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_25 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_25 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_25 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_26 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_26 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_26 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_26 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_26 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_27 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_27 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_27 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_27 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_27 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_28 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_28 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_28 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_28 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_28 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_29 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_29 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_29 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_29 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_29 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module FF_WIDTH32_30 ( clk, data_i, data_o );
  input [31:0] data_i;
  output [31:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[31]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[31]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[31]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[30]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[30]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[30]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[29]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[29]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[29]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[28]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[28]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[28]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[27]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[27]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[27]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[26]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[26]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[26]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[25]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[25]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[25]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[24]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[24]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[24]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[23]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[23]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[23]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[22]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[22]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[22]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[21]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[21]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[21]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[20]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[20]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[20]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[19]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[19]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[19]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[18]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[18]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[18]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[17]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[17]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[17]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[16]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[16]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[16]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[15]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[15]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[15]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[14]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[14]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[14]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[13]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[13]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[13]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[12]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[12]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[12]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[11]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[11]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[11]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[10]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[10]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[10]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[9]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[9]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[9]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[8]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[8]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[8]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[7]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[7]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[7]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[6]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[6]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[6]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[5]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[5]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[5]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[4]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[4]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[4]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[3]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[3]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[3]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[2]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[2]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[2]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[1]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[1]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[1]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module FF_30 ( clk, data_i, data_o );
  input [0:0] data_i;
  output [0:0] data_o;
  input clk;


  \**SEQGEN**  \data_reg[0]  ( .clear(1'b0), .preset(1'b0), .next_state(
        data_i[0]), .clocked_on(clk), .data_in(1'b0), .enable(1'b0), .Q(
        data_o[0]), .synch_clear(1'b0), .synch_preset(1'b0), .synch_toggle(
        1'b0), .synch_enable(1'b1) );
endmodule


module cam_word_30 ( clk, reset, read, dec_read_index, write, dec_write_index, 
        write_data, search, search_data, search_results, read_results, 
        read_value );
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  input clk, reset, read, dec_read_index, write, dec_write_index, search;
  output search_results, read_results;
  wire   N0, valid_i, valid_o, N1, N2, N3, N4, N5, N6, N7, N8, N9;
  wire   [31:0] data_i;

  FF_WIDTH32_30 data_ff ( .clk(clk), .data_i(data_i), .data_o(read_value) );
  FF_30 valid_ff ( .clk(clk), .data_i(valid_i), .data_o(valid_o) );
  EQ_UNS_OP eq_56_2 ( .A(search_data), .B(read_value), .Z(N1) );
  SELECT_OP C68 ( .DATA1(1'b0), .DATA2(1'b1), .DATA3(valid_o), .CONTROL1(N0), 
        .CONTROL2(N8), .CONTROL3(N6), .Z(valid_i) );
  GTECH_BUF B_0 ( .A(reset), .Z(N0) );
  SELECT_OP C69 ( .DATA1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .DATA2(write_data), .DATA3(read_value), .CONTROL1(N0), .CONTROL2(N8), 
        .CONTROL3(N6), .Z(data_i) );
  GTECH_AND2 C72 ( .A(search), .B(N1), .Z(N2) );
  GTECH_BUF B_1 ( .A(N2), .Z(search_results) );
  GTECH_AND2 C74 ( .A(N9), .B(valid_o), .Z(N3) );
  GTECH_AND2 C75 ( .A(read), .B(dec_read_index), .Z(N9) );
  GTECH_BUF B_2 ( .A(N3), .Z(read_results) );
  GTECH_AND2 C77 ( .A(dec_write_index), .B(write), .Z(N4) );
  GTECH_OR2 C80 ( .A(N4), .B(reset), .Z(N5) );
  GTECH_NOT I_0 ( .A(N5), .Z(N6) );
  GTECH_NOT I_1 ( .A(reset), .Z(N7) );
  GTECH_AND2 C83 ( .A(N4), .B(N7), .Z(N8) );
endmodule


module decoder_5_32_0 ( decoder_i, decoder_o );
  input [4:0] decoder_i;
  output [31:0] decoder_o;
  wire   N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29,
         N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43,
         N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96;

  GTECH_AND2 C4 ( .A(decoder_i[4]), .B(decoder_i[3]), .Z(N0) );
  GTECH_AND2 C5 ( .A(decoder_i[2]), .B(decoder_i[1]), .Z(N1) );
  GTECH_AND2 C6 ( .A(N0), .B(N1), .Z(N2) );
  GTECH_AND2 C7 ( .A(N2), .B(decoder_i[0]), .Z(N3) );
  GTECH_OR2 C17 ( .A(N88), .B(N89), .Z(N4) );
  GTECH_OR2 C18 ( .A(N90), .B(N91), .Z(N5) );
  GTECH_OR2 C19 ( .A(N4), .B(N5), .Z(N6) );
  GTECH_OR2 C20 ( .A(N6), .B(decoder_i[0]), .Z(N7) );
  GTECH_OR2 C32 ( .A(N90), .B(decoder_i[1]), .Z(N9) );
  GTECH_OR2 C33 ( .A(N4), .B(N9), .Z(N10) );
  GTECH_OR2 C34 ( .A(N10), .B(N92), .Z(N11) );
  GTECH_OR2 C47 ( .A(N10), .B(decoder_i[0]), .Z(N13) );
  GTECH_OR2 C59 ( .A(decoder_i[2]), .B(N91), .Z(N15) );
  GTECH_OR2 C60 ( .A(N4), .B(N15), .Z(N16) );
  GTECH_OR2 C61 ( .A(N16), .B(N92), .Z(N17) );
  GTECH_OR2 C74 ( .A(N16), .B(decoder_i[0]), .Z(N19) );
  GTECH_OR2 C85 ( .A(decoder_i[2]), .B(decoder_i[1]), .Z(N21) );
  GTECH_OR2 C86 ( .A(N4), .B(N21), .Z(N22) );
  GTECH_OR2 C87 ( .A(N22), .B(N92), .Z(N23) );
  GTECH_OR2 C99 ( .A(N22), .B(decoder_i[0]), .Z(N25) );
  GTECH_OR2 C110 ( .A(N88), .B(decoder_i[3]), .Z(N27) );
  GTECH_OR2 C112 ( .A(N27), .B(N5), .Z(N28) );
  GTECH_OR2 C113 ( .A(N28), .B(N92), .Z(N29) );
  GTECH_OR2 C126 ( .A(N28), .B(decoder_i[0]), .Z(N31) );
  GTECH_OR2 C138 ( .A(N27), .B(N9), .Z(N33) );
  GTECH_OR2 C139 ( .A(N33), .B(N92), .Z(N34) );
  GTECH_OR2 C151 ( .A(N33), .B(decoder_i[0]), .Z(N36) );
  GTECH_OR2 C163 ( .A(N27), .B(N15), .Z(N38) );
  GTECH_OR2 C164 ( .A(N38), .B(N92), .Z(N39) );
  GTECH_OR2 C176 ( .A(N38), .B(decoder_i[0]), .Z(N41) );
  GTECH_OR2 C187 ( .A(N27), .B(N21), .Z(N43) );
  GTECH_OR2 C188 ( .A(N43), .B(N92), .Z(N44) );
  GTECH_OR2 C199 ( .A(N43), .B(decoder_i[0]), .Z(N46) );
  GTECH_OR2 C210 ( .A(decoder_i[4]), .B(N89), .Z(N48) );
  GTECH_OR2 C212 ( .A(N48), .B(N5), .Z(N49) );
  GTECH_OR2 C213 ( .A(N49), .B(N92), .Z(N50) );
  GTECH_OR2 C226 ( .A(N49), .B(decoder_i[0]), .Z(N52) );
  GTECH_OR2 C238 ( .A(N48), .B(N9), .Z(N54) );
  GTECH_OR2 C239 ( .A(N54), .B(N92), .Z(N55) );
  GTECH_OR2 C251 ( .A(N54), .B(decoder_i[0]), .Z(N57) );
  GTECH_OR2 C263 ( .A(N48), .B(N15), .Z(N59) );
  GTECH_OR2 C264 ( .A(N59), .B(N92), .Z(N60) );
  GTECH_OR2 C276 ( .A(N59), .B(decoder_i[0]), .Z(N62) );
  GTECH_OR2 C287 ( .A(N48), .B(N21), .Z(N64) );
  GTECH_OR2 C288 ( .A(N64), .B(N92), .Z(N65) );
  GTECH_OR2 C299 ( .A(N64), .B(decoder_i[0]), .Z(N67) );
  GTECH_OR2 C309 ( .A(decoder_i[4]), .B(decoder_i[3]), .Z(N69) );
  GTECH_OR2 C311 ( .A(N69), .B(N5), .Z(N70) );
  GTECH_OR2 C312 ( .A(N70), .B(N92), .Z(N71) );
  GTECH_OR2 C324 ( .A(N70), .B(decoder_i[0]), .Z(N73) );
  GTECH_OR2 C335 ( .A(N69), .B(N9), .Z(N75) );
  GTECH_OR2 C336 ( .A(N75), .B(N92), .Z(N76) );
  GTECH_OR2 C347 ( .A(N75), .B(decoder_i[0]), .Z(N78) );
  GTECH_OR2 C358 ( .A(N69), .B(N15), .Z(N80) );
  GTECH_OR2 C359 ( .A(N80), .B(N92), .Z(N81) );
  GTECH_OR2 C370 ( .A(N80), .B(decoder_i[0]), .Z(N83) );
  GTECH_OR2 C380 ( .A(N69), .B(N21), .Z(N85) );
  GTECH_OR2 C381 ( .A(N85), .B(N92), .Z(N86) );
  GTECH_AND2 C393 ( .A(N88), .B(N89), .Z(N93) );
  GTECH_AND2 C394 ( .A(N90), .B(N91), .Z(N94) );
  GTECH_AND2 C395 ( .A(N93), .B(N94), .Z(N95) );
  GTECH_AND2 C396 ( .A(N95), .B(N92), .Z(N96) );
  GTECH_BUF B_0 ( .A(N3), .Z(decoder_o[31]) );
  GTECH_NOT I_0 ( .A(N7), .Z(N8) );
  GTECH_BUF B_1 ( .A(N8), .Z(decoder_o[30]) );
  GTECH_NOT I_1 ( .A(N11), .Z(N12) );
  GTECH_BUF B_2 ( .A(N12), .Z(decoder_o[29]) );
  GTECH_NOT I_2 ( .A(N13), .Z(N14) );
  GTECH_BUF B_3 ( .A(N14), .Z(decoder_o[28]) );
  GTECH_NOT I_3 ( .A(N17), .Z(N18) );
  GTECH_BUF B_4 ( .A(N18), .Z(decoder_o[27]) );
  GTECH_NOT I_4 ( .A(N19), .Z(N20) );
  GTECH_BUF B_5 ( .A(N20), .Z(decoder_o[26]) );
  GTECH_NOT I_5 ( .A(N23), .Z(N24) );
  GTECH_BUF B_6 ( .A(N24), .Z(decoder_o[25]) );
  GTECH_NOT I_6 ( .A(N25), .Z(N26) );
  GTECH_BUF B_7 ( .A(N26), .Z(decoder_o[24]) );
  GTECH_NOT I_7 ( .A(N29), .Z(N30) );
  GTECH_BUF B_8 ( .A(N30), .Z(decoder_o[23]) );
  GTECH_NOT I_8 ( .A(N31), .Z(N32) );
  GTECH_BUF B_9 ( .A(N32), .Z(decoder_o[22]) );
  GTECH_NOT I_9 ( .A(N34), .Z(N35) );
  GTECH_BUF B_10 ( .A(N35), .Z(decoder_o[21]) );
  GTECH_NOT I_10 ( .A(N36), .Z(N37) );
  GTECH_BUF B_11 ( .A(N37), .Z(decoder_o[20]) );
  GTECH_NOT I_11 ( .A(N39), .Z(N40) );
  GTECH_BUF B_12 ( .A(N40), .Z(decoder_o[19]) );
  GTECH_NOT I_12 ( .A(N41), .Z(N42) );
  GTECH_BUF B_13 ( .A(N42), .Z(decoder_o[18]) );
  GTECH_NOT I_13 ( .A(N44), .Z(N45) );
  GTECH_BUF B_14 ( .A(N45), .Z(decoder_o[17]) );
  GTECH_NOT I_14 ( .A(N46), .Z(N47) );
  GTECH_BUF B_15 ( .A(N47), .Z(decoder_o[16]) );
  GTECH_NOT I_15 ( .A(N50), .Z(N51) );
  GTECH_BUF B_16 ( .A(N51), .Z(decoder_o[15]) );
  GTECH_NOT I_16 ( .A(N52), .Z(N53) );
  GTECH_BUF B_17 ( .A(N53), .Z(decoder_o[14]) );
  GTECH_NOT I_17 ( .A(N55), .Z(N56) );
  GTECH_BUF B_18 ( .A(N56), .Z(decoder_o[13]) );
  GTECH_NOT I_18 ( .A(N57), .Z(N58) );
  GTECH_BUF B_19 ( .A(N58), .Z(decoder_o[12]) );
  GTECH_NOT I_19 ( .A(N60), .Z(N61) );
  GTECH_BUF B_20 ( .A(N61), .Z(decoder_o[11]) );
  GTECH_NOT I_20 ( .A(N62), .Z(N63) );
  GTECH_BUF B_21 ( .A(N63), .Z(decoder_o[10]) );
  GTECH_NOT I_21 ( .A(N65), .Z(N66) );
  GTECH_BUF B_22 ( .A(N66), .Z(decoder_o[9]) );
  GTECH_NOT I_22 ( .A(N67), .Z(N68) );
  GTECH_BUF B_23 ( .A(N68), .Z(decoder_o[8]) );
  GTECH_NOT I_23 ( .A(N71), .Z(N72) );
  GTECH_BUF B_24 ( .A(N72), .Z(decoder_o[7]) );
  GTECH_NOT I_24 ( .A(N73), .Z(N74) );
  GTECH_BUF B_25 ( .A(N74), .Z(decoder_o[6]) );
  GTECH_NOT I_25 ( .A(N76), .Z(N77) );
  GTECH_BUF B_26 ( .A(N77), .Z(decoder_o[5]) );
  GTECH_NOT I_26 ( .A(N78), .Z(N79) );
  GTECH_BUF B_27 ( .A(N79), .Z(decoder_o[4]) );
  GTECH_NOT I_27 ( .A(N81), .Z(N82) );
  GTECH_BUF B_28 ( .A(N82), .Z(decoder_o[3]) );
  GTECH_NOT I_28 ( .A(N83), .Z(N84) );
  GTECH_BUF B_29 ( .A(N84), .Z(decoder_o[2]) );
  GTECH_NOT I_29 ( .A(N86), .Z(N87) );
  GTECH_BUF B_30 ( .A(N87), .Z(decoder_o[1]) );
  GTECH_NOT I_30 ( .A(decoder_i[4]), .Z(N88) );
  GTECH_NOT I_31 ( .A(decoder_i[3]), .Z(N89) );
  GTECH_NOT I_32 ( .A(decoder_i[2]), .Z(N90) );
  GTECH_NOT I_33 ( .A(decoder_i[1]), .Z(N91) );
  GTECH_NOT I_34 ( .A(decoder_i[0]), .Z(N92) );
  GTECH_BUF B_31 ( .A(N96), .Z(decoder_o[0]) );
endmodule


module cam ( reset, clk, read, read_index, write, write_index, write_data, 
        search, search_data, read_valid, read_value, search_valid, 
        search_index );
  input [4:0] read_index;
  input [4:0] write_index;
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  output [4:0] search_index;
  input reset, clk, read, write, search;
  output read_valid, search_valid;
  wire   \read_value_mux[31][31] , \read_value_mux[31][30] ,
         \read_value_mux[31][29] , \read_value_mux[31][28] ,
         \read_value_mux[31][27] , \read_value_mux[31][26] ,
         \read_value_mux[31][25] , \read_value_mux[31][24] ,
         \read_value_mux[31][23] , \read_value_mux[31][22] ,
         \read_value_mux[31][21] , \read_value_mux[31][20] ,
         \read_value_mux[31][19] , \read_value_mux[31][18] ,
         \read_value_mux[31][17] , \read_value_mux[31][16] ,
         \read_value_mux[31][15] , \read_value_mux[31][14] ,
         \read_value_mux[31][13] , \read_value_mux[31][12] ,
         \read_value_mux[31][11] , \read_value_mux[31][10] ,
         \read_value_mux[31][9] , \read_value_mux[31][8] ,
         \read_value_mux[31][7] , \read_value_mux[31][6] ,
         \read_value_mux[31][5] , \read_value_mux[31][4] ,
         \read_value_mux[31][3] , \read_value_mux[31][2] ,
         \read_value_mux[31][1] , \read_value_mux[31][0] ,
         \read_value_mux[30][31] , \read_value_mux[30][30] ,
         \read_value_mux[30][29] , \read_value_mux[30][28] ,
         \read_value_mux[30][27] , \read_value_mux[30][26] ,
         \read_value_mux[30][25] , \read_value_mux[30][24] ,
         \read_value_mux[30][23] , \read_value_mux[30][22] ,
         \read_value_mux[30][21] , \read_value_mux[30][20] ,
         \read_value_mux[30][19] , \read_value_mux[30][18] ,
         \read_value_mux[30][17] , \read_value_mux[30][16] ,
         \read_value_mux[30][15] , \read_value_mux[30][14] ,
         \read_value_mux[30][13] , \read_value_mux[30][12] ,
         \read_value_mux[30][11] , \read_value_mux[30][10] ,
         \read_value_mux[30][9] , \read_value_mux[30][8] ,
         \read_value_mux[30][7] , \read_value_mux[30][6] ,
         \read_value_mux[30][5] , \read_value_mux[30][4] ,
         \read_value_mux[30][3] , \read_value_mux[30][2] ,
         \read_value_mux[30][1] , \read_value_mux[30][0] ,
         \read_value_mux[29][31] , \read_value_mux[29][30] ,
         \read_value_mux[29][29] , \read_value_mux[29][28] ,
         \read_value_mux[29][27] , \read_value_mux[29][26] ,
         \read_value_mux[29][25] , \read_value_mux[29][24] ,
         \read_value_mux[29][23] , \read_value_mux[29][22] ,
         \read_value_mux[29][21] , \read_value_mux[29][20] ,
         \read_value_mux[29][19] , \read_value_mux[29][18] ,
         \read_value_mux[29][17] , \read_value_mux[29][16] ,
         \read_value_mux[29][15] , \read_value_mux[29][14] ,
         \read_value_mux[29][13] , \read_value_mux[29][12] ,
         \read_value_mux[29][11] , \read_value_mux[29][10] ,
         \read_value_mux[29][9] , \read_value_mux[29][8] ,
         \read_value_mux[29][7] , \read_value_mux[29][6] ,
         \read_value_mux[29][5] , \read_value_mux[29][4] ,
         \read_value_mux[29][3] , \read_value_mux[29][2] ,
         \read_value_mux[29][1] , \read_value_mux[29][0] ,
         \read_value_mux[28][31] , \read_value_mux[28][30] ,
         \read_value_mux[28][29] , \read_value_mux[28][28] ,
         \read_value_mux[28][27] , \read_value_mux[28][26] ,
         \read_value_mux[28][25] , \read_value_mux[28][24] ,
         \read_value_mux[28][23] , \read_value_mux[28][22] ,
         \read_value_mux[28][21] , \read_value_mux[28][20] ,
         \read_value_mux[28][19] , \read_value_mux[28][18] ,
         \read_value_mux[28][17] , \read_value_mux[28][16] ,
         \read_value_mux[28][15] , \read_value_mux[28][14] ,
         \read_value_mux[28][13] , \read_value_mux[28][12] ,
         \read_value_mux[28][11] , \read_value_mux[28][10] ,
         \read_value_mux[28][9] , \read_value_mux[28][8] ,
         \read_value_mux[28][7] , \read_value_mux[28][6] ,
         \read_value_mux[28][5] , \read_value_mux[28][4] ,
         \read_value_mux[28][3] , \read_value_mux[28][2] ,
         \read_value_mux[28][1] , \read_value_mux[28][0] ,
         \read_value_mux[27][31] , \read_value_mux[27][30] ,
         \read_value_mux[27][29] , \read_value_mux[27][28] ,
         \read_value_mux[27][27] , \read_value_mux[27][26] ,
         \read_value_mux[27][25] , \read_value_mux[27][24] ,
         \read_value_mux[27][23] , \read_value_mux[27][22] ,
         \read_value_mux[27][21] , \read_value_mux[27][20] ,
         \read_value_mux[27][19] , \read_value_mux[27][18] ,
         \read_value_mux[27][17] , \read_value_mux[27][16] ,
         \read_value_mux[27][15] , \read_value_mux[27][14] ,
         \read_value_mux[27][13] , \read_value_mux[27][12] ,
         \read_value_mux[27][11] , \read_value_mux[27][10] ,
         \read_value_mux[27][9] , \read_value_mux[27][8] ,
         \read_value_mux[27][7] , \read_value_mux[27][6] ,
         \read_value_mux[27][5] , \read_value_mux[27][4] ,
         \read_value_mux[27][3] , \read_value_mux[27][2] ,
         \read_value_mux[27][1] , \read_value_mux[27][0] ,
         \read_value_mux[26][31] , \read_value_mux[26][30] ,
         \read_value_mux[26][29] , \read_value_mux[26][28] ,
         \read_value_mux[26][27] , \read_value_mux[26][26] ,
         \read_value_mux[26][25] , \read_value_mux[26][24] ,
         \read_value_mux[26][23] , \read_value_mux[26][22] ,
         \read_value_mux[26][21] , \read_value_mux[26][20] ,
         \read_value_mux[26][19] , \read_value_mux[26][18] ,
         \read_value_mux[26][17] , \read_value_mux[26][16] ,
         \read_value_mux[26][15] , \read_value_mux[26][14] ,
         \read_value_mux[26][13] , \read_value_mux[26][12] ,
         \read_value_mux[26][11] , \read_value_mux[26][10] ,
         \read_value_mux[26][9] , \read_value_mux[26][8] ,
         \read_value_mux[26][7] , \read_value_mux[26][6] ,
         \read_value_mux[26][5] , \read_value_mux[26][4] ,
         \read_value_mux[26][3] , \read_value_mux[26][2] ,
         \read_value_mux[26][1] , \read_value_mux[26][0] ,
         \read_value_mux[25][31] , \read_value_mux[25][30] ,
         \read_value_mux[25][29] , \read_value_mux[25][28] ,
         \read_value_mux[25][27] , \read_value_mux[25][26] ,
         \read_value_mux[25][25] , \read_value_mux[25][24] ,
         \read_value_mux[25][23] , \read_value_mux[25][22] ,
         \read_value_mux[25][21] , \read_value_mux[25][20] ,
         \read_value_mux[25][19] , \read_value_mux[25][18] ,
         \read_value_mux[25][17] , \read_value_mux[25][16] ,
         \read_value_mux[25][15] , \read_value_mux[25][14] ,
         \read_value_mux[25][13] , \read_value_mux[25][12] ,
         \read_value_mux[25][11] , \read_value_mux[25][10] ,
         \read_value_mux[25][9] , \read_value_mux[25][8] ,
         \read_value_mux[25][7] , \read_value_mux[25][6] ,
         \read_value_mux[25][5] , \read_value_mux[25][4] ,
         \read_value_mux[25][3] , \read_value_mux[25][2] ,
         \read_value_mux[25][1] , \read_value_mux[25][0] ,
         \read_value_mux[24][31] , \read_value_mux[24][30] ,
         \read_value_mux[24][29] , \read_value_mux[24][28] ,
         \read_value_mux[24][27] , \read_value_mux[24][26] ,
         \read_value_mux[24][25] , \read_value_mux[24][24] ,
         \read_value_mux[24][23] , \read_value_mux[24][22] ,
         \read_value_mux[24][21] , \read_value_mux[24][20] ,
         \read_value_mux[24][19] , \read_value_mux[24][18] ,
         \read_value_mux[24][17] , \read_value_mux[24][16] ,
         \read_value_mux[24][15] , \read_value_mux[24][14] ,
         \read_value_mux[24][13] , \read_value_mux[24][12] ,
         \read_value_mux[24][11] , \read_value_mux[24][10] ,
         \read_value_mux[24][9] , \read_value_mux[24][8] ,
         \read_value_mux[24][7] , \read_value_mux[24][6] ,
         \read_value_mux[24][5] , \read_value_mux[24][4] ,
         \read_value_mux[24][3] , \read_value_mux[24][2] ,
         \read_value_mux[24][1] , \read_value_mux[24][0] ,
         \read_value_mux[23][31] , \read_value_mux[23][30] ,
         \read_value_mux[23][29] , \read_value_mux[23][28] ,
         \read_value_mux[23][27] , \read_value_mux[23][26] ,
         \read_value_mux[23][25] , \read_value_mux[23][24] ,
         \read_value_mux[23][23] , \read_value_mux[23][22] ,
         \read_value_mux[23][21] , \read_value_mux[23][20] ,
         \read_value_mux[23][19] , \read_value_mux[23][18] ,
         \read_value_mux[23][17] , \read_value_mux[23][16] ,
         \read_value_mux[23][15] , \read_value_mux[23][14] ,
         \read_value_mux[23][13] , \read_value_mux[23][12] ,
         \read_value_mux[23][11] , \read_value_mux[23][10] ,
         \read_value_mux[23][9] , \read_value_mux[23][8] ,
         \read_value_mux[23][7] , \read_value_mux[23][6] ,
         \read_value_mux[23][5] , \read_value_mux[23][4] ,
         \read_value_mux[23][3] , \read_value_mux[23][2] ,
         \read_value_mux[23][1] , \read_value_mux[23][0] ,
         \read_value_mux[22][31] , \read_value_mux[22][30] ,
         \read_value_mux[22][29] , \read_value_mux[22][28] ,
         \read_value_mux[22][27] , \read_value_mux[22][26] ,
         \read_value_mux[22][25] , \read_value_mux[22][24] ,
         \read_value_mux[22][23] , \read_value_mux[22][22] ,
         \read_value_mux[22][21] , \read_value_mux[22][20] ,
         \read_value_mux[22][19] , \read_value_mux[22][18] ,
         \read_value_mux[22][17] , \read_value_mux[22][16] ,
         \read_value_mux[22][15] , \read_value_mux[22][14] ,
         \read_value_mux[22][13] , \read_value_mux[22][12] ,
         \read_value_mux[22][11] , \read_value_mux[22][10] ,
         \read_value_mux[22][9] , \read_value_mux[22][8] ,
         \read_value_mux[22][7] , \read_value_mux[22][6] ,
         \read_value_mux[22][5] , \read_value_mux[22][4] ,
         \read_value_mux[22][3] , \read_value_mux[22][2] ,
         \read_value_mux[22][1] , \read_value_mux[22][0] ,
         \read_value_mux[21][31] , \read_value_mux[21][30] ,
         \read_value_mux[21][29] , \read_value_mux[21][28] ,
         \read_value_mux[21][27] , \read_value_mux[21][26] ,
         \read_value_mux[21][25] , \read_value_mux[21][24] ,
         \read_value_mux[21][23] , \read_value_mux[21][22] ,
         \read_value_mux[21][21] , \read_value_mux[21][20] ,
         \read_value_mux[21][19] , \read_value_mux[21][18] ,
         \read_value_mux[21][17] , \read_value_mux[21][16] ,
         \read_value_mux[21][15] , \read_value_mux[21][14] ,
         \read_value_mux[21][13] , \read_value_mux[21][12] ,
         \read_value_mux[21][11] , \read_value_mux[21][10] ,
         \read_value_mux[21][9] , \read_value_mux[21][8] ,
         \read_value_mux[21][7] , \read_value_mux[21][6] ,
         \read_value_mux[21][5] , \read_value_mux[21][4] ,
         \read_value_mux[21][3] , \read_value_mux[21][2] ,
         \read_value_mux[21][1] , \read_value_mux[21][0] ,
         \read_value_mux[20][31] , \read_value_mux[20][30] ,
         \read_value_mux[20][29] , \read_value_mux[20][28] ,
         \read_value_mux[20][27] , \read_value_mux[20][26] ,
         \read_value_mux[20][25] , \read_value_mux[20][24] ,
         \read_value_mux[20][23] , \read_value_mux[20][22] ,
         \read_value_mux[20][21] , \read_value_mux[20][20] ,
         \read_value_mux[20][19] , \read_value_mux[20][18] ,
         \read_value_mux[20][17] , \read_value_mux[20][16] ,
         \read_value_mux[20][15] , \read_value_mux[20][14] ,
         \read_value_mux[20][13] , \read_value_mux[20][12] ,
         \read_value_mux[20][11] , \read_value_mux[20][10] ,
         \read_value_mux[20][9] , \read_value_mux[20][8] ,
         \read_value_mux[20][7] , \read_value_mux[20][6] ,
         \read_value_mux[20][5] , \read_value_mux[20][4] ,
         \read_value_mux[20][3] , \read_value_mux[20][2] ,
         \read_value_mux[20][1] , \read_value_mux[20][0] ,
         \read_value_mux[19][31] , \read_value_mux[19][30] ,
         \read_value_mux[19][29] , \read_value_mux[19][28] ,
         \read_value_mux[19][27] , \read_value_mux[19][26] ,
         \read_value_mux[19][25] , \read_value_mux[19][24] ,
         \read_value_mux[19][23] , \read_value_mux[19][22] ,
         \read_value_mux[19][21] , \read_value_mux[19][20] ,
         \read_value_mux[19][19] , \read_value_mux[19][18] ,
         \read_value_mux[19][17] , \read_value_mux[19][16] ,
         \read_value_mux[19][15] , \read_value_mux[19][14] ,
         \read_value_mux[19][13] , \read_value_mux[19][12] ,
         \read_value_mux[19][11] , \read_value_mux[19][10] ,
         \read_value_mux[19][9] , \read_value_mux[19][8] ,
         \read_value_mux[19][7] , \read_value_mux[19][6] ,
         \read_value_mux[19][5] , \read_value_mux[19][4] ,
         \read_value_mux[19][3] , \read_value_mux[19][2] ,
         \read_value_mux[19][1] , \read_value_mux[19][0] ,
         \read_value_mux[18][31] , \read_value_mux[18][30] ,
         \read_value_mux[18][29] , \read_value_mux[18][28] ,
         \read_value_mux[18][27] , \read_value_mux[18][26] ,
         \read_value_mux[18][25] , \read_value_mux[18][24] ,
         \read_value_mux[18][23] , \read_value_mux[18][22] ,
         \read_value_mux[18][21] , \read_value_mux[18][20] ,
         \read_value_mux[18][19] , \read_value_mux[18][18] ,
         \read_value_mux[18][17] , \read_value_mux[18][16] ,
         \read_value_mux[18][15] , \read_value_mux[18][14] ,
         \read_value_mux[18][13] , \read_value_mux[18][12] ,
         \read_value_mux[18][11] , \read_value_mux[18][10] ,
         \read_value_mux[18][9] , \read_value_mux[18][8] ,
         \read_value_mux[18][7] , \read_value_mux[18][6] ,
         \read_value_mux[18][5] , \read_value_mux[18][4] ,
         \read_value_mux[18][3] , \read_value_mux[18][2] ,
         \read_value_mux[18][1] , \read_value_mux[18][0] ,
         \read_value_mux[17][31] , \read_value_mux[17][30] ,
         \read_value_mux[17][29] , \read_value_mux[17][28] ,
         \read_value_mux[17][27] , \read_value_mux[17][26] ,
         \read_value_mux[17][25] , \read_value_mux[17][24] ,
         \read_value_mux[17][23] , \read_value_mux[17][22] ,
         \read_value_mux[17][21] , \read_value_mux[17][20] ,
         \read_value_mux[17][19] , \read_value_mux[17][18] ,
         \read_value_mux[17][17] , \read_value_mux[17][16] ,
         \read_value_mux[17][15] , \read_value_mux[17][14] ,
         \read_value_mux[17][13] , \read_value_mux[17][12] ,
         \read_value_mux[17][11] , \read_value_mux[17][10] ,
         \read_value_mux[17][9] , \read_value_mux[17][8] ,
         \read_value_mux[17][7] , \read_value_mux[17][6] ,
         \read_value_mux[17][5] , \read_value_mux[17][4] ,
         \read_value_mux[17][3] , \read_value_mux[17][2] ,
         \read_value_mux[17][1] , \read_value_mux[17][0] ,
         \read_value_mux[16][31] , \read_value_mux[16][30] ,
         \read_value_mux[16][29] , \read_value_mux[16][28] ,
         \read_value_mux[16][27] , \read_value_mux[16][26] ,
         \read_value_mux[16][25] , \read_value_mux[16][24] ,
         \read_value_mux[16][23] , \read_value_mux[16][22] ,
         \read_value_mux[16][21] , \read_value_mux[16][20] ,
         \read_value_mux[16][19] , \read_value_mux[16][18] ,
         \read_value_mux[16][17] , \read_value_mux[16][16] ,
         \read_value_mux[16][15] , \read_value_mux[16][14] ,
         \read_value_mux[16][13] , \read_value_mux[16][12] ,
         \read_value_mux[16][11] , \read_value_mux[16][10] ,
         \read_value_mux[16][9] , \read_value_mux[16][8] ,
         \read_value_mux[16][7] , \read_value_mux[16][6] ,
         \read_value_mux[16][5] , \read_value_mux[16][4] ,
         \read_value_mux[16][3] , \read_value_mux[16][2] ,
         \read_value_mux[16][1] , \read_value_mux[16][0] ,
         \read_value_mux[15][31] , \read_value_mux[15][30] ,
         \read_value_mux[15][29] , \read_value_mux[15][28] ,
         \read_value_mux[15][27] , \read_value_mux[15][26] ,
         \read_value_mux[15][25] , \read_value_mux[15][24] ,
         \read_value_mux[15][23] , \read_value_mux[15][22] ,
         \read_value_mux[15][21] , \read_value_mux[15][20] ,
         \read_value_mux[15][19] , \read_value_mux[15][18] ,
         \read_value_mux[15][17] , \read_value_mux[15][16] ,
         \read_value_mux[15][15] , \read_value_mux[15][14] ,
         \read_value_mux[15][13] , \read_value_mux[15][12] ,
         \read_value_mux[15][11] , \read_value_mux[15][10] ,
         \read_value_mux[15][9] , \read_value_mux[15][8] ,
         \read_value_mux[15][7] , \read_value_mux[15][6] ,
         \read_value_mux[15][5] , \read_value_mux[15][4] ,
         \read_value_mux[15][3] , \read_value_mux[15][2] ,
         \read_value_mux[15][1] , \read_value_mux[15][0] ,
         \read_value_mux[14][31] , \read_value_mux[14][30] ,
         \read_value_mux[14][29] , \read_value_mux[14][28] ,
         \read_value_mux[14][27] , \read_value_mux[14][26] ,
         \read_value_mux[14][25] , \read_value_mux[14][24] ,
         \read_value_mux[14][23] , \read_value_mux[14][22] ,
         \read_value_mux[14][21] , \read_value_mux[14][20] ,
         \read_value_mux[14][19] , \read_value_mux[14][18] ,
         \read_value_mux[14][17] , \read_value_mux[14][16] ,
         \read_value_mux[14][15] , \read_value_mux[14][14] ,
         \read_value_mux[14][13] , \read_value_mux[14][12] ,
         \read_value_mux[14][11] , \read_value_mux[14][10] ,
         \read_value_mux[14][9] , \read_value_mux[14][8] ,
         \read_value_mux[14][7] , \read_value_mux[14][6] ,
         \read_value_mux[14][5] , \read_value_mux[14][4] ,
         \read_value_mux[14][3] , \read_value_mux[14][2] ,
         \read_value_mux[14][1] , \read_value_mux[14][0] ,
         \read_value_mux[13][31] , \read_value_mux[13][30] ,
         \read_value_mux[13][29] , \read_value_mux[13][28] ,
         \read_value_mux[13][27] , \read_value_mux[13][26] ,
         \read_value_mux[13][25] , \read_value_mux[13][24] ,
         \read_value_mux[13][23] , \read_value_mux[13][22] ,
         \read_value_mux[13][21] , \read_value_mux[13][20] ,
         \read_value_mux[13][19] , \read_value_mux[13][18] ,
         \read_value_mux[13][17] , \read_value_mux[13][16] ,
         \read_value_mux[13][15] , \read_value_mux[13][14] ,
         \read_value_mux[13][13] , \read_value_mux[13][12] ,
         \read_value_mux[13][11] , \read_value_mux[13][10] ,
         \read_value_mux[13][9] , \read_value_mux[13][8] ,
         \read_value_mux[13][7] , \read_value_mux[13][6] ,
         \read_value_mux[13][5] , \read_value_mux[13][4] ,
         \read_value_mux[13][3] , \read_value_mux[13][2] ,
         \read_value_mux[13][1] , \read_value_mux[13][0] ,
         \read_value_mux[12][31] , \read_value_mux[12][30] ,
         \read_value_mux[12][29] , \read_value_mux[12][28] ,
         \read_value_mux[12][27] , \read_value_mux[12][26] ,
         \read_value_mux[12][25] , \read_value_mux[12][24] ,
         \read_value_mux[12][23] , \read_value_mux[12][22] ,
         \read_value_mux[12][21] , \read_value_mux[12][20] ,
         \read_value_mux[12][19] , \read_value_mux[12][18] ,
         \read_value_mux[12][17] , \read_value_mux[12][16] ,
         \read_value_mux[12][15] , \read_value_mux[12][14] ,
         \read_value_mux[12][13] , \read_value_mux[12][12] ,
         \read_value_mux[12][11] , \read_value_mux[12][10] ,
         \read_value_mux[12][9] , \read_value_mux[12][8] ,
         \read_value_mux[12][7] , \read_value_mux[12][6] ,
         \read_value_mux[12][5] , \read_value_mux[12][4] ,
         \read_value_mux[12][3] , \read_value_mux[12][2] ,
         \read_value_mux[12][1] , \read_value_mux[12][0] ,
         \read_value_mux[11][31] , \read_value_mux[11][30] ,
         \read_value_mux[11][29] , \read_value_mux[11][28] ,
         \read_value_mux[11][27] , \read_value_mux[11][26] ,
         \read_value_mux[11][25] , \read_value_mux[11][24] ,
         \read_value_mux[11][23] , \read_value_mux[11][22] ,
         \read_value_mux[11][21] , \read_value_mux[11][20] ,
         \read_value_mux[11][19] , \read_value_mux[11][18] ,
         \read_value_mux[11][17] , \read_value_mux[11][16] ,
         \read_value_mux[11][15] , \read_value_mux[11][14] ,
         \read_value_mux[11][13] , \read_value_mux[11][12] ,
         \read_value_mux[11][11] , \read_value_mux[11][10] ,
         \read_value_mux[11][9] , \read_value_mux[11][8] ,
         \read_value_mux[11][7] , \read_value_mux[11][6] ,
         \read_value_mux[11][5] , \read_value_mux[11][4] ,
         \read_value_mux[11][3] , \read_value_mux[11][2] ,
         \read_value_mux[11][1] , \read_value_mux[11][0] ,
         \read_value_mux[10][31] , \read_value_mux[10][30] ,
         \read_value_mux[10][29] , \read_value_mux[10][28] ,
         \read_value_mux[10][27] , \read_value_mux[10][26] ,
         \read_value_mux[10][25] , \read_value_mux[10][24] ,
         \read_value_mux[10][23] , \read_value_mux[10][22] ,
         \read_value_mux[10][21] , \read_value_mux[10][20] ,
         \read_value_mux[10][19] , \read_value_mux[10][18] ,
         \read_value_mux[10][17] , \read_value_mux[10][16] ,
         \read_value_mux[10][15] , \read_value_mux[10][14] ,
         \read_value_mux[10][13] , \read_value_mux[10][12] ,
         \read_value_mux[10][11] , \read_value_mux[10][10] ,
         \read_value_mux[10][9] , \read_value_mux[10][8] ,
         \read_value_mux[10][7] , \read_value_mux[10][6] ,
         \read_value_mux[10][5] , \read_value_mux[10][4] ,
         \read_value_mux[10][3] , \read_value_mux[10][2] ,
         \read_value_mux[10][1] , \read_value_mux[10][0] ,
         \read_value_mux[9][31] , \read_value_mux[9][30] ,
         \read_value_mux[9][29] , \read_value_mux[9][28] ,
         \read_value_mux[9][27] , \read_value_mux[9][26] ,
         \read_value_mux[9][25] , \read_value_mux[9][24] ,
         \read_value_mux[9][23] , \read_value_mux[9][22] ,
         \read_value_mux[9][21] , \read_value_mux[9][20] ,
         \read_value_mux[9][19] , \read_value_mux[9][18] ,
         \read_value_mux[9][17] , \read_value_mux[9][16] ,
         \read_value_mux[9][15] , \read_value_mux[9][14] ,
         \read_value_mux[9][13] , \read_value_mux[9][12] ,
         \read_value_mux[9][11] , \read_value_mux[9][10] ,
         \read_value_mux[9][9] , \read_value_mux[9][8] ,
         \read_value_mux[9][7] , \read_value_mux[9][6] ,
         \read_value_mux[9][5] , \read_value_mux[9][4] ,
         \read_value_mux[9][3] , \read_value_mux[9][2] ,
         \read_value_mux[9][1] , \read_value_mux[9][0] ,
         \read_value_mux[8][31] , \read_value_mux[8][30] ,
         \read_value_mux[8][29] , \read_value_mux[8][28] ,
         \read_value_mux[8][27] , \read_value_mux[8][26] ,
         \read_value_mux[8][25] , \read_value_mux[8][24] ,
         \read_value_mux[8][23] , \read_value_mux[8][22] ,
         \read_value_mux[8][21] , \read_value_mux[8][20] ,
         \read_value_mux[8][19] , \read_value_mux[8][18] ,
         \read_value_mux[8][17] , \read_value_mux[8][16] ,
         \read_value_mux[8][15] , \read_value_mux[8][14] ,
         \read_value_mux[8][13] , \read_value_mux[8][12] ,
         \read_value_mux[8][11] , \read_value_mux[8][10] ,
         \read_value_mux[8][9] , \read_value_mux[8][8] ,
         \read_value_mux[8][7] , \read_value_mux[8][6] ,
         \read_value_mux[8][5] , \read_value_mux[8][4] ,
         \read_value_mux[8][3] , \read_value_mux[8][2] ,
         \read_value_mux[8][1] , \read_value_mux[8][0] ,
         \read_value_mux[7][31] , \read_value_mux[7][30] ,
         \read_value_mux[7][29] , \read_value_mux[7][28] ,
         \read_value_mux[7][27] , \read_value_mux[7][26] ,
         \read_value_mux[7][25] , \read_value_mux[7][24] ,
         \read_value_mux[7][23] , \read_value_mux[7][22] ,
         \read_value_mux[7][21] , \read_value_mux[7][20] ,
         \read_value_mux[7][19] , \read_value_mux[7][18] ,
         \read_value_mux[7][17] , \read_value_mux[7][16] ,
         \read_value_mux[7][15] , \read_value_mux[7][14] ,
         \read_value_mux[7][13] , \read_value_mux[7][12] ,
         \read_value_mux[7][11] , \read_value_mux[7][10] ,
         \read_value_mux[7][9] , \read_value_mux[7][8] ,
         \read_value_mux[7][7] , \read_value_mux[7][6] ,
         \read_value_mux[7][5] , \read_value_mux[7][4] ,
         \read_value_mux[7][3] , \read_value_mux[7][2] ,
         \read_value_mux[7][1] , \read_value_mux[7][0] ,
         \read_value_mux[6][31] , \read_value_mux[6][30] ,
         \read_value_mux[6][29] , \read_value_mux[6][28] ,
         \read_value_mux[6][27] , \read_value_mux[6][26] ,
         \read_value_mux[6][25] , \read_value_mux[6][24] ,
         \read_value_mux[6][23] , \read_value_mux[6][22] ,
         \read_value_mux[6][21] , \read_value_mux[6][20] ,
         \read_value_mux[6][19] , \read_value_mux[6][18] ,
         \read_value_mux[6][17] , \read_value_mux[6][16] ,
         \read_value_mux[6][15] , \read_value_mux[6][14] ,
         \read_value_mux[6][13] , \read_value_mux[6][12] ,
         \read_value_mux[6][11] , \read_value_mux[6][10] ,
         \read_value_mux[6][9] , \read_value_mux[6][8] ,
         \read_value_mux[6][7] , \read_value_mux[6][6] ,
         \read_value_mux[6][5] , \read_value_mux[6][4] ,
         \read_value_mux[6][3] , \read_value_mux[6][2] ,
         \read_value_mux[6][1] , \read_value_mux[6][0] ,
         \read_value_mux[5][31] , \read_value_mux[5][30] ,
         \read_value_mux[5][29] , \read_value_mux[5][28] ,
         \read_value_mux[5][27] , \read_value_mux[5][26] ,
         \read_value_mux[5][25] , \read_value_mux[5][24] ,
         \read_value_mux[5][23] , \read_value_mux[5][22] ,
         \read_value_mux[5][21] , \read_value_mux[5][20] ,
         \read_value_mux[5][19] , \read_value_mux[5][18] ,
         \read_value_mux[5][17] , \read_value_mux[5][16] ,
         \read_value_mux[5][15] , \read_value_mux[5][14] ,
         \read_value_mux[5][13] , \read_value_mux[5][12] ,
         \read_value_mux[5][11] , \read_value_mux[5][10] ,
         \read_value_mux[5][9] , \read_value_mux[5][8] ,
         \read_value_mux[5][7] , \read_value_mux[5][6] ,
         \read_value_mux[5][5] , \read_value_mux[5][4] ,
         \read_value_mux[5][3] , \read_value_mux[5][2] ,
         \read_value_mux[5][1] , \read_value_mux[5][0] ,
         \read_value_mux[4][31] , \read_value_mux[4][30] ,
         \read_value_mux[4][29] , \read_value_mux[4][28] ,
         \read_value_mux[4][27] , \read_value_mux[4][26] ,
         \read_value_mux[4][25] , \read_value_mux[4][24] ,
         \read_value_mux[4][23] , \read_value_mux[4][22] ,
         \read_value_mux[4][21] , \read_value_mux[4][20] ,
         \read_value_mux[4][19] , \read_value_mux[4][18] ,
         \read_value_mux[4][17] , \read_value_mux[4][16] ,
         \read_value_mux[4][15] , \read_value_mux[4][14] ,
         \read_value_mux[4][13] , \read_value_mux[4][12] ,
         \read_value_mux[4][11] , \read_value_mux[4][10] ,
         \read_value_mux[4][9] , \read_value_mux[4][8] ,
         \read_value_mux[4][7] , \read_value_mux[4][6] ,
         \read_value_mux[4][5] , \read_value_mux[4][4] ,
         \read_value_mux[4][3] , \read_value_mux[4][2] ,
         \read_value_mux[4][1] , \read_value_mux[4][0] ,
         \read_value_mux[3][31] , \read_value_mux[3][30] ,
         \read_value_mux[3][29] , \read_value_mux[3][28] ,
         \read_value_mux[3][27] , \read_value_mux[3][26] ,
         \read_value_mux[3][25] , \read_value_mux[3][24] ,
         \read_value_mux[3][23] , \read_value_mux[3][22] ,
         \read_value_mux[3][21] , \read_value_mux[3][20] ,
         \read_value_mux[3][19] , \read_value_mux[3][18] ,
         \read_value_mux[3][17] , \read_value_mux[3][16] ,
         \read_value_mux[3][15] , \read_value_mux[3][14] ,
         \read_value_mux[3][13] , \read_value_mux[3][12] ,
         \read_value_mux[3][11] , \read_value_mux[3][10] ,
         \read_value_mux[3][9] , \read_value_mux[3][8] ,
         \read_value_mux[3][7] , \read_value_mux[3][6] ,
         \read_value_mux[3][5] , \read_value_mux[3][4] ,
         \read_value_mux[3][3] , \read_value_mux[3][2] ,
         \read_value_mux[3][1] , \read_value_mux[3][0] ,
         \read_value_mux[2][31] , \read_value_mux[2][30] ,
         \read_value_mux[2][29] , \read_value_mux[2][28] ,
         \read_value_mux[2][27] , \read_value_mux[2][26] ,
         \read_value_mux[2][25] , \read_value_mux[2][24] ,
         \read_value_mux[2][23] , \read_value_mux[2][22] ,
         \read_value_mux[2][21] , \read_value_mux[2][20] ,
         \read_value_mux[2][19] , \read_value_mux[2][18] ,
         \read_value_mux[2][17] , \read_value_mux[2][16] ,
         \read_value_mux[2][15] , \read_value_mux[2][14] ,
         \read_value_mux[2][13] , \read_value_mux[2][12] ,
         \read_value_mux[2][11] , \read_value_mux[2][10] ,
         \read_value_mux[2][9] , \read_value_mux[2][8] ,
         \read_value_mux[2][7] , \read_value_mux[2][6] ,
         \read_value_mux[2][5] , \read_value_mux[2][4] ,
         \read_value_mux[2][3] , \read_value_mux[2][2] ,
         \read_value_mux[2][1] , \read_value_mux[2][0] ,
         \read_value_mux[1][31] , \read_value_mux[1][30] ,
         \read_value_mux[1][29] , \read_value_mux[1][28] ,
         \read_value_mux[1][27] , \read_value_mux[1][26] ,
         \read_value_mux[1][25] , \read_value_mux[1][24] ,
         \read_value_mux[1][23] , \read_value_mux[1][22] ,
         \read_value_mux[1][21] , \read_value_mux[1][20] ,
         \read_value_mux[1][19] , \read_value_mux[1][18] ,
         \read_value_mux[1][17] , \read_value_mux[1][16] ,
         \read_value_mux[1][15] , \read_value_mux[1][14] ,
         \read_value_mux[1][13] , \read_value_mux[1][12] ,
         \read_value_mux[1][11] , \read_value_mux[1][10] ,
         \read_value_mux[1][9] , \read_value_mux[1][8] ,
         \read_value_mux[1][7] , \read_value_mux[1][6] ,
         \read_value_mux[1][5] , \read_value_mux[1][4] ,
         \read_value_mux[1][3] , \read_value_mux[1][2] ,
         \read_value_mux[1][1] , \read_value_mux[1][0] ,
         \read_value_mux[0][31] , \read_value_mux[0][30] ,
         \read_value_mux[0][29] , \read_value_mux[0][28] ,
         \read_value_mux[0][27] , \read_value_mux[0][26] ,
         \read_value_mux[0][25] , \read_value_mux[0][24] ,
         \read_value_mux[0][23] , \read_value_mux[0][22] ,
         \read_value_mux[0][21] , \read_value_mux[0][20] ,
         \read_value_mux[0][19] , \read_value_mux[0][18] ,
         \read_value_mux[0][17] , \read_value_mux[0][16] ,
         \read_value_mux[0][15] , \read_value_mux[0][14] ,
         \read_value_mux[0][13] , \read_value_mux[0][12] ,
         \read_value_mux[0][11] , \read_value_mux[0][10] ,
         \read_value_mux[0][9] , \read_value_mux[0][8] ,
         \read_value_mux[0][7] , \read_value_mux[0][6] ,
         \read_value_mux[0][5] , \read_value_mux[0][4] ,
         \read_value_mux[0][3] , \read_value_mux[0][2] ,
         \read_value_mux[0][1] , \read_value_mux[0][0] , N0, N1, N2, N3, N4,
         N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33,
         N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47,
         N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59;
  wire   [31:0] dec_read_index;
  wire   [31:0] dec_write_index;
  wire   [31:0] search_results;
  wire   [31:0] read_results;

  cam_word_0 \words[0]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[0]), .write(write), .dec_write_index(
        dec_write_index[0]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[0]), 
        .read_results(read_results[0]), .read_value({\read_value_mux[0][31] , 
        \read_value_mux[0][30] , \read_value_mux[0][29] , 
        \read_value_mux[0][28] , \read_value_mux[0][27] , 
        \read_value_mux[0][26] , \read_value_mux[0][25] , 
        \read_value_mux[0][24] , \read_value_mux[0][23] , 
        \read_value_mux[0][22] , \read_value_mux[0][21] , 
        \read_value_mux[0][20] , \read_value_mux[0][19] , 
        \read_value_mux[0][18] , \read_value_mux[0][17] , 
        \read_value_mux[0][16] , \read_value_mux[0][15] , 
        \read_value_mux[0][14] , \read_value_mux[0][13] , 
        \read_value_mux[0][12] , \read_value_mux[0][11] , 
        \read_value_mux[0][10] , \read_value_mux[0][9] , 
        \read_value_mux[0][8] , \read_value_mux[0][7] , \read_value_mux[0][6] , 
        \read_value_mux[0][5] , \read_value_mux[0][4] , \read_value_mux[0][3] , 
        \read_value_mux[0][2] , \read_value_mux[0][1] , \read_value_mux[0][0] }) );
  cam_word_1 \words[1]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[1]), .write(write), .dec_write_index(
        dec_write_index[1]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[1]), 
        .read_results(read_results[1]), .read_value({\read_value_mux[1][31] , 
        \read_value_mux[1][30] , \read_value_mux[1][29] , 
        \read_value_mux[1][28] , \read_value_mux[1][27] , 
        \read_value_mux[1][26] , \read_value_mux[1][25] , 
        \read_value_mux[1][24] , \read_value_mux[1][23] , 
        \read_value_mux[1][22] , \read_value_mux[1][21] , 
        \read_value_mux[1][20] , \read_value_mux[1][19] , 
        \read_value_mux[1][18] , \read_value_mux[1][17] , 
        \read_value_mux[1][16] , \read_value_mux[1][15] , 
        \read_value_mux[1][14] , \read_value_mux[1][13] , 
        \read_value_mux[1][12] , \read_value_mux[1][11] , 
        \read_value_mux[1][10] , \read_value_mux[1][9] , 
        \read_value_mux[1][8] , \read_value_mux[1][7] , \read_value_mux[1][6] , 
        \read_value_mux[1][5] , \read_value_mux[1][4] , \read_value_mux[1][3] , 
        \read_value_mux[1][2] , \read_value_mux[1][1] , \read_value_mux[1][0] }) );
  cam_word_2 \words[2]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[2]), .write(write), .dec_write_index(
        dec_write_index[2]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[2]), 
        .read_results(read_results[2]), .read_value({\read_value_mux[2][31] , 
        \read_value_mux[2][30] , \read_value_mux[2][29] , 
        \read_value_mux[2][28] , \read_value_mux[2][27] , 
        \read_value_mux[2][26] , \read_value_mux[2][25] , 
        \read_value_mux[2][24] , \read_value_mux[2][23] , 
        \read_value_mux[2][22] , \read_value_mux[2][21] , 
        \read_value_mux[2][20] , \read_value_mux[2][19] , 
        \read_value_mux[2][18] , \read_value_mux[2][17] , 
        \read_value_mux[2][16] , \read_value_mux[2][15] , 
        \read_value_mux[2][14] , \read_value_mux[2][13] , 
        \read_value_mux[2][12] , \read_value_mux[2][11] , 
        \read_value_mux[2][10] , \read_value_mux[2][9] , 
        \read_value_mux[2][8] , \read_value_mux[2][7] , \read_value_mux[2][6] , 
        \read_value_mux[2][5] , \read_value_mux[2][4] , \read_value_mux[2][3] , 
        \read_value_mux[2][2] , \read_value_mux[2][1] , \read_value_mux[2][0] }) );
  cam_word_3 \words[3]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[3]), .write(write), .dec_write_index(
        dec_write_index[3]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[3]), 
        .read_results(read_results[3]), .read_value({\read_value_mux[3][31] , 
        \read_value_mux[3][30] , \read_value_mux[3][29] , 
        \read_value_mux[3][28] , \read_value_mux[3][27] , 
        \read_value_mux[3][26] , \read_value_mux[3][25] , 
        \read_value_mux[3][24] , \read_value_mux[3][23] , 
        \read_value_mux[3][22] , \read_value_mux[3][21] , 
        \read_value_mux[3][20] , \read_value_mux[3][19] , 
        \read_value_mux[3][18] , \read_value_mux[3][17] , 
        \read_value_mux[3][16] , \read_value_mux[3][15] , 
        \read_value_mux[3][14] , \read_value_mux[3][13] , 
        \read_value_mux[3][12] , \read_value_mux[3][11] , 
        \read_value_mux[3][10] , \read_value_mux[3][9] , 
        \read_value_mux[3][8] , \read_value_mux[3][7] , \read_value_mux[3][6] , 
        \read_value_mux[3][5] , \read_value_mux[3][4] , \read_value_mux[3][3] , 
        \read_value_mux[3][2] , \read_value_mux[3][1] , \read_value_mux[3][0] }) );
  cam_word_4 \words[4]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[4]), .write(write), .dec_write_index(
        dec_write_index[4]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[4]), 
        .read_results(read_results[4]), .read_value({\read_value_mux[4][31] , 
        \read_value_mux[4][30] , \read_value_mux[4][29] , 
        \read_value_mux[4][28] , \read_value_mux[4][27] , 
        \read_value_mux[4][26] , \read_value_mux[4][25] , 
        \read_value_mux[4][24] , \read_value_mux[4][23] , 
        \read_value_mux[4][22] , \read_value_mux[4][21] , 
        \read_value_mux[4][20] , \read_value_mux[4][19] , 
        \read_value_mux[4][18] , \read_value_mux[4][17] , 
        \read_value_mux[4][16] , \read_value_mux[4][15] , 
        \read_value_mux[4][14] , \read_value_mux[4][13] , 
        \read_value_mux[4][12] , \read_value_mux[4][11] , 
        \read_value_mux[4][10] , \read_value_mux[4][9] , 
        \read_value_mux[4][8] , \read_value_mux[4][7] , \read_value_mux[4][6] , 
        \read_value_mux[4][5] , \read_value_mux[4][4] , \read_value_mux[4][3] , 
        \read_value_mux[4][2] , \read_value_mux[4][1] , \read_value_mux[4][0] }) );
  cam_word_5 \words[5]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[5]), .write(write), .dec_write_index(
        dec_write_index[5]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[5]), 
        .read_results(read_results[5]), .read_value({\read_value_mux[5][31] , 
        \read_value_mux[5][30] , \read_value_mux[5][29] , 
        \read_value_mux[5][28] , \read_value_mux[5][27] , 
        \read_value_mux[5][26] , \read_value_mux[5][25] , 
        \read_value_mux[5][24] , \read_value_mux[5][23] , 
        \read_value_mux[5][22] , \read_value_mux[5][21] , 
        \read_value_mux[5][20] , \read_value_mux[5][19] , 
        \read_value_mux[5][18] , \read_value_mux[5][17] , 
        \read_value_mux[5][16] , \read_value_mux[5][15] , 
        \read_value_mux[5][14] , \read_value_mux[5][13] , 
        \read_value_mux[5][12] , \read_value_mux[5][11] , 
        \read_value_mux[5][10] , \read_value_mux[5][9] , 
        \read_value_mux[5][8] , \read_value_mux[5][7] , \read_value_mux[5][6] , 
        \read_value_mux[5][5] , \read_value_mux[5][4] , \read_value_mux[5][3] , 
        \read_value_mux[5][2] , \read_value_mux[5][1] , \read_value_mux[5][0] }) );
  cam_word_6 \words[6]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[6]), .write(write), .dec_write_index(
        dec_write_index[6]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[6]), 
        .read_results(read_results[6]), .read_value({\read_value_mux[6][31] , 
        \read_value_mux[6][30] , \read_value_mux[6][29] , 
        \read_value_mux[6][28] , \read_value_mux[6][27] , 
        \read_value_mux[6][26] , \read_value_mux[6][25] , 
        \read_value_mux[6][24] , \read_value_mux[6][23] , 
        \read_value_mux[6][22] , \read_value_mux[6][21] , 
        \read_value_mux[6][20] , \read_value_mux[6][19] , 
        \read_value_mux[6][18] , \read_value_mux[6][17] , 
        \read_value_mux[6][16] , \read_value_mux[6][15] , 
        \read_value_mux[6][14] , \read_value_mux[6][13] , 
        \read_value_mux[6][12] , \read_value_mux[6][11] , 
        \read_value_mux[6][10] , \read_value_mux[6][9] , 
        \read_value_mux[6][8] , \read_value_mux[6][7] , \read_value_mux[6][6] , 
        \read_value_mux[6][5] , \read_value_mux[6][4] , \read_value_mux[6][3] , 
        \read_value_mux[6][2] , \read_value_mux[6][1] , \read_value_mux[6][0] }) );
  cam_word_7 \words[7]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[7]), .write(write), .dec_write_index(
        dec_write_index[7]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[7]), 
        .read_results(read_results[7]), .read_value({\read_value_mux[7][31] , 
        \read_value_mux[7][30] , \read_value_mux[7][29] , 
        \read_value_mux[7][28] , \read_value_mux[7][27] , 
        \read_value_mux[7][26] , \read_value_mux[7][25] , 
        \read_value_mux[7][24] , \read_value_mux[7][23] , 
        \read_value_mux[7][22] , \read_value_mux[7][21] , 
        \read_value_mux[7][20] , \read_value_mux[7][19] , 
        \read_value_mux[7][18] , \read_value_mux[7][17] , 
        \read_value_mux[7][16] , \read_value_mux[7][15] , 
        \read_value_mux[7][14] , \read_value_mux[7][13] , 
        \read_value_mux[7][12] , \read_value_mux[7][11] , 
        \read_value_mux[7][10] , \read_value_mux[7][9] , 
        \read_value_mux[7][8] , \read_value_mux[7][7] , \read_value_mux[7][6] , 
        \read_value_mux[7][5] , \read_value_mux[7][4] , \read_value_mux[7][3] , 
        \read_value_mux[7][2] , \read_value_mux[7][1] , \read_value_mux[7][0] }) );
  cam_word_8 \words[8]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[8]), .write(write), .dec_write_index(
        dec_write_index[8]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[8]), 
        .read_results(read_results[8]), .read_value({\read_value_mux[8][31] , 
        \read_value_mux[8][30] , \read_value_mux[8][29] , 
        \read_value_mux[8][28] , \read_value_mux[8][27] , 
        \read_value_mux[8][26] , \read_value_mux[8][25] , 
        \read_value_mux[8][24] , \read_value_mux[8][23] , 
        \read_value_mux[8][22] , \read_value_mux[8][21] , 
        \read_value_mux[8][20] , \read_value_mux[8][19] , 
        \read_value_mux[8][18] , \read_value_mux[8][17] , 
        \read_value_mux[8][16] , \read_value_mux[8][15] , 
        \read_value_mux[8][14] , \read_value_mux[8][13] , 
        \read_value_mux[8][12] , \read_value_mux[8][11] , 
        \read_value_mux[8][10] , \read_value_mux[8][9] , 
        \read_value_mux[8][8] , \read_value_mux[8][7] , \read_value_mux[8][6] , 
        \read_value_mux[8][5] , \read_value_mux[8][4] , \read_value_mux[8][3] , 
        \read_value_mux[8][2] , \read_value_mux[8][1] , \read_value_mux[8][0] }) );
  cam_word_9 \words[9]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[9]), .write(write), .dec_write_index(
        dec_write_index[9]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[9]), 
        .read_results(read_results[9]), .read_value({\read_value_mux[9][31] , 
        \read_value_mux[9][30] , \read_value_mux[9][29] , 
        \read_value_mux[9][28] , \read_value_mux[9][27] , 
        \read_value_mux[9][26] , \read_value_mux[9][25] , 
        \read_value_mux[9][24] , \read_value_mux[9][23] , 
        \read_value_mux[9][22] , \read_value_mux[9][21] , 
        \read_value_mux[9][20] , \read_value_mux[9][19] , 
        \read_value_mux[9][18] , \read_value_mux[9][17] , 
        \read_value_mux[9][16] , \read_value_mux[9][15] , 
        \read_value_mux[9][14] , \read_value_mux[9][13] , 
        \read_value_mux[9][12] , \read_value_mux[9][11] , 
        \read_value_mux[9][10] , \read_value_mux[9][9] , 
        \read_value_mux[9][8] , \read_value_mux[9][7] , \read_value_mux[9][6] , 
        \read_value_mux[9][5] , \read_value_mux[9][4] , \read_value_mux[9][3] , 
        \read_value_mux[9][2] , \read_value_mux[9][1] , \read_value_mux[9][0] }) );
  cam_word_10 \words[10]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[10]), .write(write), .dec_write_index(
        dec_write_index[10]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[10]), 
        .read_results(read_results[10]), .read_value({\read_value_mux[10][31] , 
        \read_value_mux[10][30] , \read_value_mux[10][29] , 
        \read_value_mux[10][28] , \read_value_mux[10][27] , 
        \read_value_mux[10][26] , \read_value_mux[10][25] , 
        \read_value_mux[10][24] , \read_value_mux[10][23] , 
        \read_value_mux[10][22] , \read_value_mux[10][21] , 
        \read_value_mux[10][20] , \read_value_mux[10][19] , 
        \read_value_mux[10][18] , \read_value_mux[10][17] , 
        \read_value_mux[10][16] , \read_value_mux[10][15] , 
        \read_value_mux[10][14] , \read_value_mux[10][13] , 
        \read_value_mux[10][12] , \read_value_mux[10][11] , 
        \read_value_mux[10][10] , \read_value_mux[10][9] , 
        \read_value_mux[10][8] , \read_value_mux[10][7] , 
        \read_value_mux[10][6] , \read_value_mux[10][5] , 
        \read_value_mux[10][4] , \read_value_mux[10][3] , 
        \read_value_mux[10][2] , \read_value_mux[10][1] , 
        \read_value_mux[10][0] }) );
  cam_word_11 \words[11]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[11]), .write(write), .dec_write_index(
        dec_write_index[11]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[11]), 
        .read_results(read_results[11]), .read_value({\read_value_mux[11][31] , 
        \read_value_mux[11][30] , \read_value_mux[11][29] , 
        \read_value_mux[11][28] , \read_value_mux[11][27] , 
        \read_value_mux[11][26] , \read_value_mux[11][25] , 
        \read_value_mux[11][24] , \read_value_mux[11][23] , 
        \read_value_mux[11][22] , \read_value_mux[11][21] , 
        \read_value_mux[11][20] , \read_value_mux[11][19] , 
        \read_value_mux[11][18] , \read_value_mux[11][17] , 
        \read_value_mux[11][16] , \read_value_mux[11][15] , 
        \read_value_mux[11][14] , \read_value_mux[11][13] , 
        \read_value_mux[11][12] , \read_value_mux[11][11] , 
        \read_value_mux[11][10] , \read_value_mux[11][9] , 
        \read_value_mux[11][8] , \read_value_mux[11][7] , 
        \read_value_mux[11][6] , \read_value_mux[11][5] , 
        \read_value_mux[11][4] , \read_value_mux[11][3] , 
        \read_value_mux[11][2] , \read_value_mux[11][1] , 
        \read_value_mux[11][0] }) );
  cam_word_12 \words[12]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[12]), .write(write), .dec_write_index(
        dec_write_index[12]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[12]), 
        .read_results(read_results[12]), .read_value({\read_value_mux[12][31] , 
        \read_value_mux[12][30] , \read_value_mux[12][29] , 
        \read_value_mux[12][28] , \read_value_mux[12][27] , 
        \read_value_mux[12][26] , \read_value_mux[12][25] , 
        \read_value_mux[12][24] , \read_value_mux[12][23] , 
        \read_value_mux[12][22] , \read_value_mux[12][21] , 
        \read_value_mux[12][20] , \read_value_mux[12][19] , 
        \read_value_mux[12][18] , \read_value_mux[12][17] , 
        \read_value_mux[12][16] , \read_value_mux[12][15] , 
        \read_value_mux[12][14] , \read_value_mux[12][13] , 
        \read_value_mux[12][12] , \read_value_mux[12][11] , 
        \read_value_mux[12][10] , \read_value_mux[12][9] , 
        \read_value_mux[12][8] , \read_value_mux[12][7] , 
        \read_value_mux[12][6] , \read_value_mux[12][5] , 
        \read_value_mux[12][4] , \read_value_mux[12][3] , 
        \read_value_mux[12][2] , \read_value_mux[12][1] , 
        \read_value_mux[12][0] }) );
  cam_word_13 \words[13]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[13]), .write(write), .dec_write_index(
        dec_write_index[13]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[13]), 
        .read_results(read_results[13]), .read_value({\read_value_mux[13][31] , 
        \read_value_mux[13][30] , \read_value_mux[13][29] , 
        \read_value_mux[13][28] , \read_value_mux[13][27] , 
        \read_value_mux[13][26] , \read_value_mux[13][25] , 
        \read_value_mux[13][24] , \read_value_mux[13][23] , 
        \read_value_mux[13][22] , \read_value_mux[13][21] , 
        \read_value_mux[13][20] , \read_value_mux[13][19] , 
        \read_value_mux[13][18] , \read_value_mux[13][17] , 
        \read_value_mux[13][16] , \read_value_mux[13][15] , 
        \read_value_mux[13][14] , \read_value_mux[13][13] , 
        \read_value_mux[13][12] , \read_value_mux[13][11] , 
        \read_value_mux[13][10] , \read_value_mux[13][9] , 
        \read_value_mux[13][8] , \read_value_mux[13][7] , 
        \read_value_mux[13][6] , \read_value_mux[13][5] , 
        \read_value_mux[13][4] , \read_value_mux[13][3] , 
        \read_value_mux[13][2] , \read_value_mux[13][1] , 
        \read_value_mux[13][0] }) );
  cam_word_14 \words[14]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[14]), .write(write), .dec_write_index(
        dec_write_index[14]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[14]), 
        .read_results(read_results[14]), .read_value({\read_value_mux[14][31] , 
        \read_value_mux[14][30] , \read_value_mux[14][29] , 
        \read_value_mux[14][28] , \read_value_mux[14][27] , 
        \read_value_mux[14][26] , \read_value_mux[14][25] , 
        \read_value_mux[14][24] , \read_value_mux[14][23] , 
        \read_value_mux[14][22] , \read_value_mux[14][21] , 
        \read_value_mux[14][20] , \read_value_mux[14][19] , 
        \read_value_mux[14][18] , \read_value_mux[14][17] , 
        \read_value_mux[14][16] , \read_value_mux[14][15] , 
        \read_value_mux[14][14] , \read_value_mux[14][13] , 
        \read_value_mux[14][12] , \read_value_mux[14][11] , 
        \read_value_mux[14][10] , \read_value_mux[14][9] , 
        \read_value_mux[14][8] , \read_value_mux[14][7] , 
        \read_value_mux[14][6] , \read_value_mux[14][5] , 
        \read_value_mux[14][4] , \read_value_mux[14][3] , 
        \read_value_mux[14][2] , \read_value_mux[14][1] , 
        \read_value_mux[14][0] }) );
  cam_word_15 \words[15]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[15]), .write(write), .dec_write_index(
        dec_write_index[15]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[15]), 
        .read_results(read_results[15]), .read_value({\read_value_mux[15][31] , 
        \read_value_mux[15][30] , \read_value_mux[15][29] , 
        \read_value_mux[15][28] , \read_value_mux[15][27] , 
        \read_value_mux[15][26] , \read_value_mux[15][25] , 
        \read_value_mux[15][24] , \read_value_mux[15][23] , 
        \read_value_mux[15][22] , \read_value_mux[15][21] , 
        \read_value_mux[15][20] , \read_value_mux[15][19] , 
        \read_value_mux[15][18] , \read_value_mux[15][17] , 
        \read_value_mux[15][16] , \read_value_mux[15][15] , 
        \read_value_mux[15][14] , \read_value_mux[15][13] , 
        \read_value_mux[15][12] , \read_value_mux[15][11] , 
        \read_value_mux[15][10] , \read_value_mux[15][9] , 
        \read_value_mux[15][8] , \read_value_mux[15][7] , 
        \read_value_mux[15][6] , \read_value_mux[15][5] , 
        \read_value_mux[15][4] , \read_value_mux[15][3] , 
        \read_value_mux[15][2] , \read_value_mux[15][1] , 
        \read_value_mux[15][0] }) );
  cam_word_16 \words[16]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[16]), .write(write), .dec_write_index(
        dec_write_index[16]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[16]), 
        .read_results(read_results[16]), .read_value({\read_value_mux[16][31] , 
        \read_value_mux[16][30] , \read_value_mux[16][29] , 
        \read_value_mux[16][28] , \read_value_mux[16][27] , 
        \read_value_mux[16][26] , \read_value_mux[16][25] , 
        \read_value_mux[16][24] , \read_value_mux[16][23] , 
        \read_value_mux[16][22] , \read_value_mux[16][21] , 
        \read_value_mux[16][20] , \read_value_mux[16][19] , 
        \read_value_mux[16][18] , \read_value_mux[16][17] , 
        \read_value_mux[16][16] , \read_value_mux[16][15] , 
        \read_value_mux[16][14] , \read_value_mux[16][13] , 
        \read_value_mux[16][12] , \read_value_mux[16][11] , 
        \read_value_mux[16][10] , \read_value_mux[16][9] , 
        \read_value_mux[16][8] , \read_value_mux[16][7] , 
        \read_value_mux[16][6] , \read_value_mux[16][5] , 
        \read_value_mux[16][4] , \read_value_mux[16][3] , 
        \read_value_mux[16][2] , \read_value_mux[16][1] , 
        \read_value_mux[16][0] }) );
  cam_word_17 \words[17]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[17]), .write(write), .dec_write_index(
        dec_write_index[17]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[17]), 
        .read_results(read_results[17]), .read_value({\read_value_mux[17][31] , 
        \read_value_mux[17][30] , \read_value_mux[17][29] , 
        \read_value_mux[17][28] , \read_value_mux[17][27] , 
        \read_value_mux[17][26] , \read_value_mux[17][25] , 
        \read_value_mux[17][24] , \read_value_mux[17][23] , 
        \read_value_mux[17][22] , \read_value_mux[17][21] , 
        \read_value_mux[17][20] , \read_value_mux[17][19] , 
        \read_value_mux[17][18] , \read_value_mux[17][17] , 
        \read_value_mux[17][16] , \read_value_mux[17][15] , 
        \read_value_mux[17][14] , \read_value_mux[17][13] , 
        \read_value_mux[17][12] , \read_value_mux[17][11] , 
        \read_value_mux[17][10] , \read_value_mux[17][9] , 
        \read_value_mux[17][8] , \read_value_mux[17][7] , 
        \read_value_mux[17][6] , \read_value_mux[17][5] , 
        \read_value_mux[17][4] , \read_value_mux[17][3] , 
        \read_value_mux[17][2] , \read_value_mux[17][1] , 
        \read_value_mux[17][0] }) );
  cam_word_18 \words[18]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[18]), .write(write), .dec_write_index(
        dec_write_index[18]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[18]), 
        .read_results(read_results[18]), .read_value({\read_value_mux[18][31] , 
        \read_value_mux[18][30] , \read_value_mux[18][29] , 
        \read_value_mux[18][28] , \read_value_mux[18][27] , 
        \read_value_mux[18][26] , \read_value_mux[18][25] , 
        \read_value_mux[18][24] , \read_value_mux[18][23] , 
        \read_value_mux[18][22] , \read_value_mux[18][21] , 
        \read_value_mux[18][20] , \read_value_mux[18][19] , 
        \read_value_mux[18][18] , \read_value_mux[18][17] , 
        \read_value_mux[18][16] , \read_value_mux[18][15] , 
        \read_value_mux[18][14] , \read_value_mux[18][13] , 
        \read_value_mux[18][12] , \read_value_mux[18][11] , 
        \read_value_mux[18][10] , \read_value_mux[18][9] , 
        \read_value_mux[18][8] , \read_value_mux[18][7] , 
        \read_value_mux[18][6] , \read_value_mux[18][5] , 
        \read_value_mux[18][4] , \read_value_mux[18][3] , 
        \read_value_mux[18][2] , \read_value_mux[18][1] , 
        \read_value_mux[18][0] }) );
  cam_word_19 \words[19]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[19]), .write(write), .dec_write_index(
        dec_write_index[19]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[19]), 
        .read_results(read_results[19]), .read_value({\read_value_mux[19][31] , 
        \read_value_mux[19][30] , \read_value_mux[19][29] , 
        \read_value_mux[19][28] , \read_value_mux[19][27] , 
        \read_value_mux[19][26] , \read_value_mux[19][25] , 
        \read_value_mux[19][24] , \read_value_mux[19][23] , 
        \read_value_mux[19][22] , \read_value_mux[19][21] , 
        \read_value_mux[19][20] , \read_value_mux[19][19] , 
        \read_value_mux[19][18] , \read_value_mux[19][17] , 
        \read_value_mux[19][16] , \read_value_mux[19][15] , 
        \read_value_mux[19][14] , \read_value_mux[19][13] , 
        \read_value_mux[19][12] , \read_value_mux[19][11] , 
        \read_value_mux[19][10] , \read_value_mux[19][9] , 
        \read_value_mux[19][8] , \read_value_mux[19][7] , 
        \read_value_mux[19][6] , \read_value_mux[19][5] , 
        \read_value_mux[19][4] , \read_value_mux[19][3] , 
        \read_value_mux[19][2] , \read_value_mux[19][1] , 
        \read_value_mux[19][0] }) );
  cam_word_20 \words[20]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[20]), .write(write), .dec_write_index(
        dec_write_index[20]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[20]), 
        .read_results(read_results[20]), .read_value({\read_value_mux[20][31] , 
        \read_value_mux[20][30] , \read_value_mux[20][29] , 
        \read_value_mux[20][28] , \read_value_mux[20][27] , 
        \read_value_mux[20][26] , \read_value_mux[20][25] , 
        \read_value_mux[20][24] , \read_value_mux[20][23] , 
        \read_value_mux[20][22] , \read_value_mux[20][21] , 
        \read_value_mux[20][20] , \read_value_mux[20][19] , 
        \read_value_mux[20][18] , \read_value_mux[20][17] , 
        \read_value_mux[20][16] , \read_value_mux[20][15] , 
        \read_value_mux[20][14] , \read_value_mux[20][13] , 
        \read_value_mux[20][12] , \read_value_mux[20][11] , 
        \read_value_mux[20][10] , \read_value_mux[20][9] , 
        \read_value_mux[20][8] , \read_value_mux[20][7] , 
        \read_value_mux[20][6] , \read_value_mux[20][5] , 
        \read_value_mux[20][4] , \read_value_mux[20][3] , 
        \read_value_mux[20][2] , \read_value_mux[20][1] , 
        \read_value_mux[20][0] }) );
  cam_word_21 \words[21]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[21]), .write(write), .dec_write_index(
        dec_write_index[21]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[21]), 
        .read_results(read_results[21]), .read_value({\read_value_mux[21][31] , 
        \read_value_mux[21][30] , \read_value_mux[21][29] , 
        \read_value_mux[21][28] , \read_value_mux[21][27] , 
        \read_value_mux[21][26] , \read_value_mux[21][25] , 
        \read_value_mux[21][24] , \read_value_mux[21][23] , 
        \read_value_mux[21][22] , \read_value_mux[21][21] , 
        \read_value_mux[21][20] , \read_value_mux[21][19] , 
        \read_value_mux[21][18] , \read_value_mux[21][17] , 
        \read_value_mux[21][16] , \read_value_mux[21][15] , 
        \read_value_mux[21][14] , \read_value_mux[21][13] , 
        \read_value_mux[21][12] , \read_value_mux[21][11] , 
        \read_value_mux[21][10] , \read_value_mux[21][9] , 
        \read_value_mux[21][8] , \read_value_mux[21][7] , 
        \read_value_mux[21][6] , \read_value_mux[21][5] , 
        \read_value_mux[21][4] , \read_value_mux[21][3] , 
        \read_value_mux[21][2] , \read_value_mux[21][1] , 
        \read_value_mux[21][0] }) );
  cam_word_22 \words[22]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[22]), .write(write), .dec_write_index(
        dec_write_index[22]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[22]), 
        .read_results(read_results[22]), .read_value({\read_value_mux[22][31] , 
        \read_value_mux[22][30] , \read_value_mux[22][29] , 
        \read_value_mux[22][28] , \read_value_mux[22][27] , 
        \read_value_mux[22][26] , \read_value_mux[22][25] , 
        \read_value_mux[22][24] , \read_value_mux[22][23] , 
        \read_value_mux[22][22] , \read_value_mux[22][21] , 
        \read_value_mux[22][20] , \read_value_mux[22][19] , 
        \read_value_mux[22][18] , \read_value_mux[22][17] , 
        \read_value_mux[22][16] , \read_value_mux[22][15] , 
        \read_value_mux[22][14] , \read_value_mux[22][13] , 
        \read_value_mux[22][12] , \read_value_mux[22][11] , 
        \read_value_mux[22][10] , \read_value_mux[22][9] , 
        \read_value_mux[22][8] , \read_value_mux[22][7] , 
        \read_value_mux[22][6] , \read_value_mux[22][5] , 
        \read_value_mux[22][4] , \read_value_mux[22][3] , 
        \read_value_mux[22][2] , \read_value_mux[22][1] , 
        \read_value_mux[22][0] }) );
  cam_word_23 \words[23]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[23]), .write(write), .dec_write_index(
        dec_write_index[23]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[23]), 
        .read_results(read_results[23]), .read_value({\read_value_mux[23][31] , 
        \read_value_mux[23][30] , \read_value_mux[23][29] , 
        \read_value_mux[23][28] , \read_value_mux[23][27] , 
        \read_value_mux[23][26] , \read_value_mux[23][25] , 
        \read_value_mux[23][24] , \read_value_mux[23][23] , 
        \read_value_mux[23][22] , \read_value_mux[23][21] , 
        \read_value_mux[23][20] , \read_value_mux[23][19] , 
        \read_value_mux[23][18] , \read_value_mux[23][17] , 
        \read_value_mux[23][16] , \read_value_mux[23][15] , 
        \read_value_mux[23][14] , \read_value_mux[23][13] , 
        \read_value_mux[23][12] , \read_value_mux[23][11] , 
        \read_value_mux[23][10] , \read_value_mux[23][9] , 
        \read_value_mux[23][8] , \read_value_mux[23][7] , 
        \read_value_mux[23][6] , \read_value_mux[23][5] , 
        \read_value_mux[23][4] , \read_value_mux[23][3] , 
        \read_value_mux[23][2] , \read_value_mux[23][1] , 
        \read_value_mux[23][0] }) );
  cam_word_24 \words[24]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[24]), .write(write), .dec_write_index(
        dec_write_index[24]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[24]), 
        .read_results(read_results[24]), .read_value({\read_value_mux[24][31] , 
        \read_value_mux[24][30] , \read_value_mux[24][29] , 
        \read_value_mux[24][28] , \read_value_mux[24][27] , 
        \read_value_mux[24][26] , \read_value_mux[24][25] , 
        \read_value_mux[24][24] , \read_value_mux[24][23] , 
        \read_value_mux[24][22] , \read_value_mux[24][21] , 
        \read_value_mux[24][20] , \read_value_mux[24][19] , 
        \read_value_mux[24][18] , \read_value_mux[24][17] , 
        \read_value_mux[24][16] , \read_value_mux[24][15] , 
        \read_value_mux[24][14] , \read_value_mux[24][13] , 
        \read_value_mux[24][12] , \read_value_mux[24][11] , 
        \read_value_mux[24][10] , \read_value_mux[24][9] , 
        \read_value_mux[24][8] , \read_value_mux[24][7] , 
        \read_value_mux[24][6] , \read_value_mux[24][5] , 
        \read_value_mux[24][4] , \read_value_mux[24][3] , 
        \read_value_mux[24][2] , \read_value_mux[24][1] , 
        \read_value_mux[24][0] }) );
  cam_word_25 \words[25]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[25]), .write(write), .dec_write_index(
        dec_write_index[25]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[25]), 
        .read_results(read_results[25]), .read_value({\read_value_mux[25][31] , 
        \read_value_mux[25][30] , \read_value_mux[25][29] , 
        \read_value_mux[25][28] , \read_value_mux[25][27] , 
        \read_value_mux[25][26] , \read_value_mux[25][25] , 
        \read_value_mux[25][24] , \read_value_mux[25][23] , 
        \read_value_mux[25][22] , \read_value_mux[25][21] , 
        \read_value_mux[25][20] , \read_value_mux[25][19] , 
        \read_value_mux[25][18] , \read_value_mux[25][17] , 
        \read_value_mux[25][16] , \read_value_mux[25][15] , 
        \read_value_mux[25][14] , \read_value_mux[25][13] , 
        \read_value_mux[25][12] , \read_value_mux[25][11] , 
        \read_value_mux[25][10] , \read_value_mux[25][9] , 
        \read_value_mux[25][8] , \read_value_mux[25][7] , 
        \read_value_mux[25][6] , \read_value_mux[25][5] , 
        \read_value_mux[25][4] , \read_value_mux[25][3] , 
        \read_value_mux[25][2] , \read_value_mux[25][1] , 
        \read_value_mux[25][0] }) );
  cam_word_26 \words[26]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[26]), .write(write), .dec_write_index(
        dec_write_index[26]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[26]), 
        .read_results(read_results[26]), .read_value({\read_value_mux[26][31] , 
        \read_value_mux[26][30] , \read_value_mux[26][29] , 
        \read_value_mux[26][28] , \read_value_mux[26][27] , 
        \read_value_mux[26][26] , \read_value_mux[26][25] , 
        \read_value_mux[26][24] , \read_value_mux[26][23] , 
        \read_value_mux[26][22] , \read_value_mux[26][21] , 
        \read_value_mux[26][20] , \read_value_mux[26][19] , 
        \read_value_mux[26][18] , \read_value_mux[26][17] , 
        \read_value_mux[26][16] , \read_value_mux[26][15] , 
        \read_value_mux[26][14] , \read_value_mux[26][13] , 
        \read_value_mux[26][12] , \read_value_mux[26][11] , 
        \read_value_mux[26][10] , \read_value_mux[26][9] , 
        \read_value_mux[26][8] , \read_value_mux[26][7] , 
        \read_value_mux[26][6] , \read_value_mux[26][5] , 
        \read_value_mux[26][4] , \read_value_mux[26][3] , 
        \read_value_mux[26][2] , \read_value_mux[26][1] , 
        \read_value_mux[26][0] }) );
  cam_word_27 \words[27]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[27]), .write(write), .dec_write_index(
        dec_write_index[27]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[27]), 
        .read_results(read_results[27]), .read_value({\read_value_mux[27][31] , 
        \read_value_mux[27][30] , \read_value_mux[27][29] , 
        \read_value_mux[27][28] , \read_value_mux[27][27] , 
        \read_value_mux[27][26] , \read_value_mux[27][25] , 
        \read_value_mux[27][24] , \read_value_mux[27][23] , 
        \read_value_mux[27][22] , \read_value_mux[27][21] , 
        \read_value_mux[27][20] , \read_value_mux[27][19] , 
        \read_value_mux[27][18] , \read_value_mux[27][17] , 
        \read_value_mux[27][16] , \read_value_mux[27][15] , 
        \read_value_mux[27][14] , \read_value_mux[27][13] , 
        \read_value_mux[27][12] , \read_value_mux[27][11] , 
        \read_value_mux[27][10] , \read_value_mux[27][9] , 
        \read_value_mux[27][8] , \read_value_mux[27][7] , 
        \read_value_mux[27][6] , \read_value_mux[27][5] , 
        \read_value_mux[27][4] , \read_value_mux[27][3] , 
        \read_value_mux[27][2] , \read_value_mux[27][1] , 
        \read_value_mux[27][0] }) );
  cam_word_28 \words[28]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[28]), .write(write), .dec_write_index(
        dec_write_index[28]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[28]), 
        .read_results(read_results[28]), .read_value({\read_value_mux[28][31] , 
        \read_value_mux[28][30] , \read_value_mux[28][29] , 
        \read_value_mux[28][28] , \read_value_mux[28][27] , 
        \read_value_mux[28][26] , \read_value_mux[28][25] , 
        \read_value_mux[28][24] , \read_value_mux[28][23] , 
        \read_value_mux[28][22] , \read_value_mux[28][21] , 
        \read_value_mux[28][20] , \read_value_mux[28][19] , 
        \read_value_mux[28][18] , \read_value_mux[28][17] , 
        \read_value_mux[28][16] , \read_value_mux[28][15] , 
        \read_value_mux[28][14] , \read_value_mux[28][13] , 
        \read_value_mux[28][12] , \read_value_mux[28][11] , 
        \read_value_mux[28][10] , \read_value_mux[28][9] , 
        \read_value_mux[28][8] , \read_value_mux[28][7] , 
        \read_value_mux[28][6] , \read_value_mux[28][5] , 
        \read_value_mux[28][4] , \read_value_mux[28][3] , 
        \read_value_mux[28][2] , \read_value_mux[28][1] , 
        \read_value_mux[28][0] }) );
  cam_word_29 \words[29]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[29]), .write(write), .dec_write_index(
        dec_write_index[29]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[29]), 
        .read_results(read_results[29]), .read_value({\read_value_mux[29][31] , 
        \read_value_mux[29][30] , \read_value_mux[29][29] , 
        \read_value_mux[29][28] , \read_value_mux[29][27] , 
        \read_value_mux[29][26] , \read_value_mux[29][25] , 
        \read_value_mux[29][24] , \read_value_mux[29][23] , 
        \read_value_mux[29][22] , \read_value_mux[29][21] , 
        \read_value_mux[29][20] , \read_value_mux[29][19] , 
        \read_value_mux[29][18] , \read_value_mux[29][17] , 
        \read_value_mux[29][16] , \read_value_mux[29][15] , 
        \read_value_mux[29][14] , \read_value_mux[29][13] , 
        \read_value_mux[29][12] , \read_value_mux[29][11] , 
        \read_value_mux[29][10] , \read_value_mux[29][9] , 
        \read_value_mux[29][8] , \read_value_mux[29][7] , 
        \read_value_mux[29][6] , \read_value_mux[29][5] , 
        \read_value_mux[29][4] , \read_value_mux[29][3] , 
        \read_value_mux[29][2] , \read_value_mux[29][1] , 
        \read_value_mux[29][0] }) );
  cam_word_30 \words[30]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[30]), .write(write), .dec_write_index(
        dec_write_index[30]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[30]), 
        .read_results(read_results[30]), .read_value({\read_value_mux[30][31] , 
        \read_value_mux[30][30] , \read_value_mux[30][29] , 
        \read_value_mux[30][28] , \read_value_mux[30][27] , 
        \read_value_mux[30][26] , \read_value_mux[30][25] , 
        \read_value_mux[30][24] , \read_value_mux[30][23] , 
        \read_value_mux[30][22] , \read_value_mux[30][21] , 
        \read_value_mux[30][20] , \read_value_mux[30][19] , 
        \read_value_mux[30][18] , \read_value_mux[30][17] , 
        \read_value_mux[30][16] , \read_value_mux[30][15] , 
        \read_value_mux[30][14] , \read_value_mux[30][13] , 
        \read_value_mux[30][12] , \read_value_mux[30][11] , 
        \read_value_mux[30][10] , \read_value_mux[30][9] , 
        \read_value_mux[30][8] , \read_value_mux[30][7] , 
        \read_value_mux[30][6] , \read_value_mux[30][5] , 
        \read_value_mux[30][4] , \read_value_mux[30][3] , 
        \read_value_mux[30][2] , \read_value_mux[30][1] , 
        \read_value_mux[30][0] }) );
  cam_word_31 \words[31]  ( .clk(clk), .reset(reset), .read(read), 
        .dec_read_index(dec_read_index[31]), .write(write), .dec_write_index(
        dec_write_index[31]), .write_data(write_data), .search(search), 
        .search_data(search_data), .search_results(search_results[31]), 
        .read_results(read_results[31]), .read_value({\read_value_mux[31][31] , 
        \read_value_mux[31][30] , \read_value_mux[31][29] , 
        \read_value_mux[31][28] , \read_value_mux[31][27] , 
        \read_value_mux[31][26] , \read_value_mux[31][25] , 
        \read_value_mux[31][24] , \read_value_mux[31][23] , 
        \read_value_mux[31][22] , \read_value_mux[31][21] , 
        \read_value_mux[31][20] , \read_value_mux[31][19] , 
        \read_value_mux[31][18] , \read_value_mux[31][17] , 
        \read_value_mux[31][16] , \read_value_mux[31][15] , 
        \read_value_mux[31][14] , \read_value_mux[31][13] , 
        \read_value_mux[31][12] , \read_value_mux[31][11] , 
        \read_value_mux[31][10] , \read_value_mux[31][9] , 
        \read_value_mux[31][8] , \read_value_mux[31][7] , 
        \read_value_mux[31][6] , \read_value_mux[31][5] , 
        \read_value_mux[31][4] , \read_value_mux[31][3] , 
        \read_value_mux[31][2] , \read_value_mux[31][1] , 
        \read_value_mux[31][0] }) );
  decoder_5_32_1 read_dcdr ( .decoder_i(read_index), .decoder_o(dec_read_index) );
  decoder_5_32_0 write_dcdr ( .decoder_i(write_index), .decoder_o(
        dec_write_index) );
  priority_encoder search_ecdr ( .inp_i(search_results), .out_o(search_index), 
        .valid_o(search_valid) );
  mux read_mux ( .data_i({\read_value_mux[31][31] , \read_value_mux[31][30] , 
        \read_value_mux[31][29] , \read_value_mux[31][28] , 
        \read_value_mux[31][27] , \read_value_mux[31][26] , 
        \read_value_mux[31][25] , \read_value_mux[31][24] , 
        \read_value_mux[31][23] , \read_value_mux[31][22] , 
        \read_value_mux[31][21] , \read_value_mux[31][20] , 
        \read_value_mux[31][19] , \read_value_mux[31][18] , 
        \read_value_mux[31][17] , \read_value_mux[31][16] , 
        \read_value_mux[31][15] , \read_value_mux[31][14] , 
        \read_value_mux[31][13] , \read_value_mux[31][12] , 
        \read_value_mux[31][11] , \read_value_mux[31][10] , 
        \read_value_mux[31][9] , \read_value_mux[31][8] , 
        \read_value_mux[31][7] , \read_value_mux[31][6] , 
        \read_value_mux[31][5] , \read_value_mux[31][4] , 
        \read_value_mux[31][3] , \read_value_mux[31][2] , 
        \read_value_mux[31][1] , \read_value_mux[31][0] , 
        \read_value_mux[30][31] , \read_value_mux[30][30] , 
        \read_value_mux[30][29] , \read_value_mux[30][28] , 
        \read_value_mux[30][27] , \read_value_mux[30][26] , 
        \read_value_mux[30][25] , \read_value_mux[30][24] , 
        \read_value_mux[30][23] , \read_value_mux[30][22] , 
        \read_value_mux[30][21] , \read_value_mux[30][20] , 
        \read_value_mux[30][19] , \read_value_mux[30][18] , 
        \read_value_mux[30][17] , \read_value_mux[30][16] , 
        \read_value_mux[30][15] , \read_value_mux[30][14] , 
        \read_value_mux[30][13] , \read_value_mux[30][12] , 
        \read_value_mux[30][11] , \read_value_mux[30][10] , 
        \read_value_mux[30][9] , \read_value_mux[30][8] , 
        \read_value_mux[30][7] , \read_value_mux[30][6] , 
        \read_value_mux[30][5] , \read_value_mux[30][4] , 
        \read_value_mux[30][3] , \read_value_mux[30][2] , 
        \read_value_mux[30][1] , \read_value_mux[30][0] , 
        \read_value_mux[29][31] , \read_value_mux[29][30] , 
        \read_value_mux[29][29] , \read_value_mux[29][28] , 
        \read_value_mux[29][27] , \read_value_mux[29][26] , 
        \read_value_mux[29][25] , \read_value_mux[29][24] , 
        \read_value_mux[29][23] , \read_value_mux[29][22] , 
        \read_value_mux[29][21] , \read_value_mux[29][20] , 
        \read_value_mux[29][19] , \read_value_mux[29][18] , 
        \read_value_mux[29][17] , \read_value_mux[29][16] , 
        \read_value_mux[29][15] , \read_value_mux[29][14] , 
        \read_value_mux[29][13] , \read_value_mux[29][12] , 
        \read_value_mux[29][11] , \read_value_mux[29][10] , 
        \read_value_mux[29][9] , \read_value_mux[29][8] , 
        \read_value_mux[29][7] , \read_value_mux[29][6] , 
        \read_value_mux[29][5] , \read_value_mux[29][4] , 
        \read_value_mux[29][3] , \read_value_mux[29][2] , 
        \read_value_mux[29][1] , \read_value_mux[29][0] , 
        \read_value_mux[28][31] , \read_value_mux[28][30] , 
        \read_value_mux[28][29] , \read_value_mux[28][28] , 
        \read_value_mux[28][27] , \read_value_mux[28][26] , 
        \read_value_mux[28][25] , \read_value_mux[28][24] , 
        \read_value_mux[28][23] , \read_value_mux[28][22] , 
        \read_value_mux[28][21] , \read_value_mux[28][20] , 
        \read_value_mux[28][19] , \read_value_mux[28][18] , 
        \read_value_mux[28][17] , \read_value_mux[28][16] , 
        \read_value_mux[28][15] , \read_value_mux[28][14] , 
        \read_value_mux[28][13] , \read_value_mux[28][12] , 
        \read_value_mux[28][11] , \read_value_mux[28][10] , 
        \read_value_mux[28][9] , \read_value_mux[28][8] , 
        \read_value_mux[28][7] , \read_value_mux[28][6] , 
        \read_value_mux[28][5] , \read_value_mux[28][4] , 
        \read_value_mux[28][3] , \read_value_mux[28][2] , 
        \read_value_mux[28][1] , \read_value_mux[28][0] , 
        \read_value_mux[27][31] , \read_value_mux[27][30] , 
        \read_value_mux[27][29] , \read_value_mux[27][28] , 
        \read_value_mux[27][27] , \read_value_mux[27][26] , 
        \read_value_mux[27][25] , \read_value_mux[27][24] , 
        \read_value_mux[27][23] , \read_value_mux[27][22] , 
        \read_value_mux[27][21] , \read_value_mux[27][20] , 
        \read_value_mux[27][19] , \read_value_mux[27][18] , 
        \read_value_mux[27][17] , \read_value_mux[27][16] , 
        \read_value_mux[27][15] , \read_value_mux[27][14] , 
        \read_value_mux[27][13] , \read_value_mux[27][12] , 
        \read_value_mux[27][11] , \read_value_mux[27][10] , 
        \read_value_mux[27][9] , \read_value_mux[27][8] , 
        \read_value_mux[27][7] , \read_value_mux[27][6] , 
        \read_value_mux[27][5] , \read_value_mux[27][4] , 
        \read_value_mux[27][3] , \read_value_mux[27][2] , 
        \read_value_mux[27][1] , \read_value_mux[27][0] , 
        \read_value_mux[26][31] , \read_value_mux[26][30] , 
        \read_value_mux[26][29] , \read_value_mux[26][28] , 
        \read_value_mux[26][27] , \read_value_mux[26][26] , 
        \read_value_mux[26][25] , \read_value_mux[26][24] , 
        \read_value_mux[26][23] , \read_value_mux[26][22] , 
        \read_value_mux[26][21] , \read_value_mux[26][20] , 
        \read_value_mux[26][19] , \read_value_mux[26][18] , 
        \read_value_mux[26][17] , \read_value_mux[26][16] , 
        \read_value_mux[26][15] , \read_value_mux[26][14] , 
        \read_value_mux[26][13] , \read_value_mux[26][12] , 
        \read_value_mux[26][11] , \read_value_mux[26][10] , 
        \read_value_mux[26][9] , \read_value_mux[26][8] , 
        \read_value_mux[26][7] , \read_value_mux[26][6] , 
        \read_value_mux[26][5] , \read_value_mux[26][4] , 
        \read_value_mux[26][3] , \read_value_mux[26][2] , 
        \read_value_mux[26][1] , \read_value_mux[26][0] , 
        \read_value_mux[25][31] , \read_value_mux[25][30] , 
        \read_value_mux[25][29] , \read_value_mux[25][28] , 
        \read_value_mux[25][27] , \read_value_mux[25][26] , 
        \read_value_mux[25][25] , \read_value_mux[25][24] , 
        \read_value_mux[25][23] , \read_value_mux[25][22] , 
        \read_value_mux[25][21] , \read_value_mux[25][20] , 
        \read_value_mux[25][19] , \read_value_mux[25][18] , 
        \read_value_mux[25][17] , \read_value_mux[25][16] , 
        \read_value_mux[25][15] , \read_value_mux[25][14] , 
        \read_value_mux[25][13] , \read_value_mux[25][12] , 
        \read_value_mux[25][11] , \read_value_mux[25][10] , 
        \read_value_mux[25][9] , \read_value_mux[25][8] , 
        \read_value_mux[25][7] , \read_value_mux[25][6] , 
        \read_value_mux[25][5] , \read_value_mux[25][4] , 
        \read_value_mux[25][3] , \read_value_mux[25][2] , 
        \read_value_mux[25][1] , \read_value_mux[25][0] , 
        \read_value_mux[24][31] , \read_value_mux[24][30] , 
        \read_value_mux[24][29] , \read_value_mux[24][28] , 
        \read_value_mux[24][27] , \read_value_mux[24][26] , 
        \read_value_mux[24][25] , \read_value_mux[24][24] , 
        \read_value_mux[24][23] , \read_value_mux[24][22] , 
        \read_value_mux[24][21] , \read_value_mux[24][20] , 
        \read_value_mux[24][19] , \read_value_mux[24][18] , 
        \read_value_mux[24][17] , \read_value_mux[24][16] , 
        \read_value_mux[24][15] , \read_value_mux[24][14] , 
        \read_value_mux[24][13] , \read_value_mux[24][12] , 
        \read_value_mux[24][11] , \read_value_mux[24][10] , 
        \read_value_mux[24][9] , \read_value_mux[24][8] , 
        \read_value_mux[24][7] , \read_value_mux[24][6] , 
        \read_value_mux[24][5] , \read_value_mux[24][4] , 
        \read_value_mux[24][3] , \read_value_mux[24][2] , 
        \read_value_mux[24][1] , \read_value_mux[24][0] , 
        \read_value_mux[23][31] , \read_value_mux[23][30] , 
        \read_value_mux[23][29] , \read_value_mux[23][28] , 
        \read_value_mux[23][27] , \read_value_mux[23][26] , 
        \read_value_mux[23][25] , \read_value_mux[23][24] , 
        \read_value_mux[23][23] , \read_value_mux[23][22] , 
        \read_value_mux[23][21] , \read_value_mux[23][20] , 
        \read_value_mux[23][19] , \read_value_mux[23][18] , 
        \read_value_mux[23][17] , \read_value_mux[23][16] , 
        \read_value_mux[23][15] , \read_value_mux[23][14] , 
        \read_value_mux[23][13] , \read_value_mux[23][12] , 
        \read_value_mux[23][11] , \read_value_mux[23][10] , 
        \read_value_mux[23][9] , \read_value_mux[23][8] , 
        \read_value_mux[23][7] , \read_value_mux[23][6] , 
        \read_value_mux[23][5] , \read_value_mux[23][4] , 
        \read_value_mux[23][3] , \read_value_mux[23][2] , 
        \read_value_mux[23][1] , \read_value_mux[23][0] , 
        \read_value_mux[22][31] , \read_value_mux[22][30] , 
        \read_value_mux[22][29] , \read_value_mux[22][28] , 
        \read_value_mux[22][27] , \read_value_mux[22][26] , 
        \read_value_mux[22][25] , \read_value_mux[22][24] , 
        \read_value_mux[22][23] , \read_value_mux[22][22] , 
        \read_value_mux[22][21] , \read_value_mux[22][20] , 
        \read_value_mux[22][19] , \read_value_mux[22][18] , 
        \read_value_mux[22][17] , \read_value_mux[22][16] , 
        \read_value_mux[22][15] , \read_value_mux[22][14] , 
        \read_value_mux[22][13] , \read_value_mux[22][12] , 
        \read_value_mux[22][11] , \read_value_mux[22][10] , 
        \read_value_mux[22][9] , \read_value_mux[22][8] , 
        \read_value_mux[22][7] , \read_value_mux[22][6] , 
        \read_value_mux[22][5] , \read_value_mux[22][4] , 
        \read_value_mux[22][3] , \read_value_mux[22][2] , 
        \read_value_mux[22][1] , \read_value_mux[22][0] , 
        \read_value_mux[21][31] , \read_value_mux[21][30] , 
        \read_value_mux[21][29] , \read_value_mux[21][28] , 
        \read_value_mux[21][27] , \read_value_mux[21][26] , 
        \read_value_mux[21][25] , \read_value_mux[21][24] , 
        \read_value_mux[21][23] , \read_value_mux[21][22] , 
        \read_value_mux[21][21] , \read_value_mux[21][20] , 
        \read_value_mux[21][19] , \read_value_mux[21][18] , 
        \read_value_mux[21][17] , \read_value_mux[21][16] , 
        \read_value_mux[21][15] , \read_value_mux[21][14] , 
        \read_value_mux[21][13] , \read_value_mux[21][12] , 
        \read_value_mux[21][11] , \read_value_mux[21][10] , 
        \read_value_mux[21][9] , \read_value_mux[21][8] , 
        \read_value_mux[21][7] , \read_value_mux[21][6] , 
        \read_value_mux[21][5] , \read_value_mux[21][4] , 
        \read_value_mux[21][3] , \read_value_mux[21][2] , 
        \read_value_mux[21][1] , \read_value_mux[21][0] , 
        \read_value_mux[20][31] , \read_value_mux[20][30] , 
        \read_value_mux[20][29] , \read_value_mux[20][28] , 
        \read_value_mux[20][27] , \read_value_mux[20][26] , 
        \read_value_mux[20][25] , \read_value_mux[20][24] , 
        \read_value_mux[20][23] , \read_value_mux[20][22] , 
        \read_value_mux[20][21] , \read_value_mux[20][20] , 
        \read_value_mux[20][19] , \read_value_mux[20][18] , 
        \read_value_mux[20][17] , \read_value_mux[20][16] , 
        \read_value_mux[20][15] , \read_value_mux[20][14] , 
        \read_value_mux[20][13] , \read_value_mux[20][12] , 
        \read_value_mux[20][11] , \read_value_mux[20][10] , 
        \read_value_mux[20][9] , \read_value_mux[20][8] , 
        \read_value_mux[20][7] , \read_value_mux[20][6] , 
        \read_value_mux[20][5] , \read_value_mux[20][4] , 
        \read_value_mux[20][3] , \read_value_mux[20][2] , 
        \read_value_mux[20][1] , \read_value_mux[20][0] , 
        \read_value_mux[19][31] , \read_value_mux[19][30] , 
        \read_value_mux[19][29] , \read_value_mux[19][28] , 
        \read_value_mux[19][27] , \read_value_mux[19][26] , 
        \read_value_mux[19][25] , \read_value_mux[19][24] , 
        \read_value_mux[19][23] , \read_value_mux[19][22] , 
        \read_value_mux[19][21] , \read_value_mux[19][20] , 
        \read_value_mux[19][19] , \read_value_mux[19][18] , 
        \read_value_mux[19][17] , \read_value_mux[19][16] , 
        \read_value_mux[19][15] , \read_value_mux[19][14] , 
        \read_value_mux[19][13] , \read_value_mux[19][12] , 
        \read_value_mux[19][11] , \read_value_mux[19][10] , 
        \read_value_mux[19][9] , \read_value_mux[19][8] , 
        \read_value_mux[19][7] , \read_value_mux[19][6] , 
        \read_value_mux[19][5] , \read_value_mux[19][4] , 
        \read_value_mux[19][3] , \read_value_mux[19][2] , 
        \read_value_mux[19][1] , \read_value_mux[19][0] , 
        \read_value_mux[18][31] , \read_value_mux[18][30] , 
        \read_value_mux[18][29] , \read_value_mux[18][28] , 
        \read_value_mux[18][27] , \read_value_mux[18][26] , 
        \read_value_mux[18][25] , \read_value_mux[18][24] , 
        \read_value_mux[18][23] , \read_value_mux[18][22] , 
        \read_value_mux[18][21] , \read_value_mux[18][20] , 
        \read_value_mux[18][19] , \read_value_mux[18][18] , 
        \read_value_mux[18][17] , \read_value_mux[18][16] , 
        \read_value_mux[18][15] , \read_value_mux[18][14] , 
        \read_value_mux[18][13] , \read_value_mux[18][12] , 
        \read_value_mux[18][11] , \read_value_mux[18][10] , 
        \read_value_mux[18][9] , \read_value_mux[18][8] , 
        \read_value_mux[18][7] , \read_value_mux[18][6] , 
        \read_value_mux[18][5] , \read_value_mux[18][4] , 
        \read_value_mux[18][3] , \read_value_mux[18][2] , 
        \read_value_mux[18][1] , \read_value_mux[18][0] , 
        \read_value_mux[17][31] , \read_value_mux[17][30] , 
        \read_value_mux[17][29] , \read_value_mux[17][28] , 
        \read_value_mux[17][27] , \read_value_mux[17][26] , 
        \read_value_mux[17][25] , \read_value_mux[17][24] , 
        \read_value_mux[17][23] , \read_value_mux[17][22] , 
        \read_value_mux[17][21] , \read_value_mux[17][20] , 
        \read_value_mux[17][19] , \read_value_mux[17][18] , 
        \read_value_mux[17][17] , \read_value_mux[17][16] , 
        \read_value_mux[17][15] , \read_value_mux[17][14] , 
        \read_value_mux[17][13] , \read_value_mux[17][12] , 
        \read_value_mux[17][11] , \read_value_mux[17][10] , 
        \read_value_mux[17][9] , \read_value_mux[17][8] , 
        \read_value_mux[17][7] , \read_value_mux[17][6] , 
        \read_value_mux[17][5] , \read_value_mux[17][4] , 
        \read_value_mux[17][3] , \read_value_mux[17][2] , 
        \read_value_mux[17][1] , \read_value_mux[17][0] , 
        \read_value_mux[16][31] , \read_value_mux[16][30] , 
        \read_value_mux[16][29] , \read_value_mux[16][28] , 
        \read_value_mux[16][27] , \read_value_mux[16][26] , 
        \read_value_mux[16][25] , \read_value_mux[16][24] , 
        \read_value_mux[16][23] , \read_value_mux[16][22] , 
        \read_value_mux[16][21] , \read_value_mux[16][20] , 
        \read_value_mux[16][19] , \read_value_mux[16][18] , 
        \read_value_mux[16][17] , \read_value_mux[16][16] , 
        \read_value_mux[16][15] , \read_value_mux[16][14] , 
        \read_value_mux[16][13] , \read_value_mux[16][12] , 
        \read_value_mux[16][11] , \read_value_mux[16][10] , 
        \read_value_mux[16][9] , \read_value_mux[16][8] , 
        \read_value_mux[16][7] , \read_value_mux[16][6] , 
        \read_value_mux[16][5] , \read_value_mux[16][4] , 
        \read_value_mux[16][3] , \read_value_mux[16][2] , 
        \read_value_mux[16][1] , \read_value_mux[16][0] , 
        \read_value_mux[15][31] , \read_value_mux[15][30] , 
        \read_value_mux[15][29] , \read_value_mux[15][28] , 
        \read_value_mux[15][27] , \read_value_mux[15][26] , 
        \read_value_mux[15][25] , \read_value_mux[15][24] , 
        \read_value_mux[15][23] , \read_value_mux[15][22] , 
        \read_value_mux[15][21] , \read_value_mux[15][20] , 
        \read_value_mux[15][19] , \read_value_mux[15][18] , 
        \read_value_mux[15][17] , \read_value_mux[15][16] , 
        \read_value_mux[15][15] , \read_value_mux[15][14] , 
        \read_value_mux[15][13] , \read_value_mux[15][12] , 
        \read_value_mux[15][11] , \read_value_mux[15][10] , 
        \read_value_mux[15][9] , \read_value_mux[15][8] , 
        \read_value_mux[15][7] , \read_value_mux[15][6] , 
        \read_value_mux[15][5] , \read_value_mux[15][4] , 
        \read_value_mux[15][3] , \read_value_mux[15][2] , 
        \read_value_mux[15][1] , \read_value_mux[15][0] , 
        \read_value_mux[14][31] , \read_value_mux[14][30] , 
        \read_value_mux[14][29] , \read_value_mux[14][28] , 
        \read_value_mux[14][27] , \read_value_mux[14][26] , 
        \read_value_mux[14][25] , \read_value_mux[14][24] , 
        \read_value_mux[14][23] , \read_value_mux[14][22] , 
        \read_value_mux[14][21] , \read_value_mux[14][20] , 
        \read_value_mux[14][19] , \read_value_mux[14][18] , 
        \read_value_mux[14][17] , \read_value_mux[14][16] , 
        \read_value_mux[14][15] , \read_value_mux[14][14] , 
        \read_value_mux[14][13] , \read_value_mux[14][12] , 
        \read_value_mux[14][11] , \read_value_mux[14][10] , 
        \read_value_mux[14][9] , \read_value_mux[14][8] , 
        \read_value_mux[14][7] , \read_value_mux[14][6] , 
        \read_value_mux[14][5] , \read_value_mux[14][4] , 
        \read_value_mux[14][3] , \read_value_mux[14][2] , 
        \read_value_mux[14][1] , \read_value_mux[14][0] , 
        \read_value_mux[13][31] , \read_value_mux[13][30] , 
        \read_value_mux[13][29] , \read_value_mux[13][28] , 
        \read_value_mux[13][27] , \read_value_mux[13][26] , 
        \read_value_mux[13][25] , \read_value_mux[13][24] , 
        \read_value_mux[13][23] , \read_value_mux[13][22] , 
        \read_value_mux[13][21] , \read_value_mux[13][20] , 
        \read_value_mux[13][19] , \read_value_mux[13][18] , 
        \read_value_mux[13][17] , \read_value_mux[13][16] , 
        \read_value_mux[13][15] , \read_value_mux[13][14] , 
        \read_value_mux[13][13] , \read_value_mux[13][12] , 
        \read_value_mux[13][11] , \read_value_mux[13][10] , 
        \read_value_mux[13][9] , \read_value_mux[13][8] , 
        \read_value_mux[13][7] , \read_value_mux[13][6] , 
        \read_value_mux[13][5] , \read_value_mux[13][4] , 
        \read_value_mux[13][3] , \read_value_mux[13][2] , 
        \read_value_mux[13][1] , \read_value_mux[13][0] , 
        \read_value_mux[12][31] , \read_value_mux[12][30] , 
        \read_value_mux[12][29] , \read_value_mux[12][28] , 
        \read_value_mux[12][27] , \read_value_mux[12][26] , 
        \read_value_mux[12][25] , \read_value_mux[12][24] , 
        \read_value_mux[12][23] , \read_value_mux[12][22] , 
        \read_value_mux[12][21] , \read_value_mux[12][20] , 
        \read_value_mux[12][19] , \read_value_mux[12][18] , 
        \read_value_mux[12][17] , \read_value_mux[12][16] , 
        \read_value_mux[12][15] , \read_value_mux[12][14] , 
        \read_value_mux[12][13] , \read_value_mux[12][12] , 
        \read_value_mux[12][11] , \read_value_mux[12][10] , 
        \read_value_mux[12][9] , \read_value_mux[12][8] , 
        \read_value_mux[12][7] , \read_value_mux[12][6] , 
        \read_value_mux[12][5] , \read_value_mux[12][4] , 
        \read_value_mux[12][3] , \read_value_mux[12][2] , 
        \read_value_mux[12][1] , \read_value_mux[12][0] , 
        \read_value_mux[11][31] , \read_value_mux[11][30] , 
        \read_value_mux[11][29] , \read_value_mux[11][28] , 
        \read_value_mux[11][27] , \read_value_mux[11][26] , 
        \read_value_mux[11][25] , \read_value_mux[11][24] , 
        \read_value_mux[11][23] , \read_value_mux[11][22] , 
        \read_value_mux[11][21] , \read_value_mux[11][20] , 
        \read_value_mux[11][19] , \read_value_mux[11][18] , 
        \read_value_mux[11][17] , \read_value_mux[11][16] , 
        \read_value_mux[11][15] , \read_value_mux[11][14] , 
        \read_value_mux[11][13] , \read_value_mux[11][12] , 
        \read_value_mux[11][11] , \read_value_mux[11][10] , 
        \read_value_mux[11][9] , \read_value_mux[11][8] , 
        \read_value_mux[11][7] , \read_value_mux[11][6] , 
        \read_value_mux[11][5] , \read_value_mux[11][4] , 
        \read_value_mux[11][3] , \read_value_mux[11][2] , 
        \read_value_mux[11][1] , \read_value_mux[11][0] , 
        \read_value_mux[10][31] , \read_value_mux[10][30] , 
        \read_value_mux[10][29] , \read_value_mux[10][28] , 
        \read_value_mux[10][27] , \read_value_mux[10][26] , 
        \read_value_mux[10][25] , \read_value_mux[10][24] , 
        \read_value_mux[10][23] , \read_value_mux[10][22] , 
        \read_value_mux[10][21] , \read_value_mux[10][20] , 
        \read_value_mux[10][19] , \read_value_mux[10][18] , 
        \read_value_mux[10][17] , \read_value_mux[10][16] , 
        \read_value_mux[10][15] , \read_value_mux[10][14] , 
        \read_value_mux[10][13] , \read_value_mux[10][12] , 
        \read_value_mux[10][11] , \read_value_mux[10][10] , 
        \read_value_mux[10][9] , \read_value_mux[10][8] , 
        \read_value_mux[10][7] , \read_value_mux[10][6] , 
        \read_value_mux[10][5] , \read_value_mux[10][4] , 
        \read_value_mux[10][3] , \read_value_mux[10][2] , 
        \read_value_mux[10][1] , \read_value_mux[10][0] , 
        \read_value_mux[9][31] , \read_value_mux[9][30] , 
        \read_value_mux[9][29] , \read_value_mux[9][28] , 
        \read_value_mux[9][27] , \read_value_mux[9][26] , 
        \read_value_mux[9][25] , \read_value_mux[9][24] , 
        \read_value_mux[9][23] , \read_value_mux[9][22] , 
        \read_value_mux[9][21] , \read_value_mux[9][20] , 
        \read_value_mux[9][19] , \read_value_mux[9][18] , 
        \read_value_mux[9][17] , \read_value_mux[9][16] , 
        \read_value_mux[9][15] , \read_value_mux[9][14] , 
        \read_value_mux[9][13] , \read_value_mux[9][12] , 
        \read_value_mux[9][11] , \read_value_mux[9][10] , 
        \read_value_mux[9][9] , \read_value_mux[9][8] , \read_value_mux[9][7] , 
        \read_value_mux[9][6] , \read_value_mux[9][5] , \read_value_mux[9][4] , 
        \read_value_mux[9][3] , \read_value_mux[9][2] , \read_value_mux[9][1] , 
        \read_value_mux[9][0] , \read_value_mux[8][31] , 
        \read_value_mux[8][30] , \read_value_mux[8][29] , 
        \read_value_mux[8][28] , \read_value_mux[8][27] , 
        \read_value_mux[8][26] , \read_value_mux[8][25] , 
        \read_value_mux[8][24] , \read_value_mux[8][23] , 
        \read_value_mux[8][22] , \read_value_mux[8][21] , 
        \read_value_mux[8][20] , \read_value_mux[8][19] , 
        \read_value_mux[8][18] , \read_value_mux[8][17] , 
        \read_value_mux[8][16] , \read_value_mux[8][15] , 
        \read_value_mux[8][14] , \read_value_mux[8][13] , 
        \read_value_mux[8][12] , \read_value_mux[8][11] , 
        \read_value_mux[8][10] , \read_value_mux[8][9] , 
        \read_value_mux[8][8] , \read_value_mux[8][7] , \read_value_mux[8][6] , 
        \read_value_mux[8][5] , \read_value_mux[8][4] , \read_value_mux[8][3] , 
        \read_value_mux[8][2] , \read_value_mux[8][1] , \read_value_mux[8][0] , 
        \read_value_mux[7][31] , \read_value_mux[7][30] , 
        \read_value_mux[7][29] , \read_value_mux[7][28] , 
        \read_value_mux[7][27] , \read_value_mux[7][26] , 
        \read_value_mux[7][25] , \read_value_mux[7][24] , 
        \read_value_mux[7][23] , \read_value_mux[7][22] , 
        \read_value_mux[7][21] , \read_value_mux[7][20] , 
        \read_value_mux[7][19] , \read_value_mux[7][18] , 
        \read_value_mux[7][17] , \read_value_mux[7][16] , 
        \read_value_mux[7][15] , \read_value_mux[7][14] , 
        \read_value_mux[7][13] , \read_value_mux[7][12] , 
        \read_value_mux[7][11] , \read_value_mux[7][10] , 
        \read_value_mux[7][9] , \read_value_mux[7][8] , \read_value_mux[7][7] , 
        \read_value_mux[7][6] , \read_value_mux[7][5] , \read_value_mux[7][4] , 
        \read_value_mux[7][3] , \read_value_mux[7][2] , \read_value_mux[7][1] , 
        \read_value_mux[7][0] , \read_value_mux[6][31] , 
        \read_value_mux[6][30] , \read_value_mux[6][29] , 
        \read_value_mux[6][28] , \read_value_mux[6][27] , 
        \read_value_mux[6][26] , \read_value_mux[6][25] , 
        \read_value_mux[6][24] , \read_value_mux[6][23] , 
        \read_value_mux[6][22] , \read_value_mux[6][21] , 
        \read_value_mux[6][20] , \read_value_mux[6][19] , 
        \read_value_mux[6][18] , \read_value_mux[6][17] , 
        \read_value_mux[6][16] , \read_value_mux[6][15] , 
        \read_value_mux[6][14] , \read_value_mux[6][13] , 
        \read_value_mux[6][12] , \read_value_mux[6][11] , 
        \read_value_mux[6][10] , \read_value_mux[6][9] , 
        \read_value_mux[6][8] , \read_value_mux[6][7] , \read_value_mux[6][6] , 
        \read_value_mux[6][5] , \read_value_mux[6][4] , \read_value_mux[6][3] , 
        \read_value_mux[6][2] , \read_value_mux[6][1] , \read_value_mux[6][0] , 
        \read_value_mux[5][31] , \read_value_mux[5][30] , 
        \read_value_mux[5][29] , \read_value_mux[5][28] , 
        \read_value_mux[5][27] , \read_value_mux[5][26] , 
        \read_value_mux[5][25] , \read_value_mux[5][24] , 
        \read_value_mux[5][23] , \read_value_mux[5][22] , 
        \read_value_mux[5][21] , \read_value_mux[5][20] , 
        \read_value_mux[5][19] , \read_value_mux[5][18] , 
        \read_value_mux[5][17] , \read_value_mux[5][16] , 
        \read_value_mux[5][15] , \read_value_mux[5][14] , 
        \read_value_mux[5][13] , \read_value_mux[5][12] , 
        \read_value_mux[5][11] , \read_value_mux[5][10] , 
        \read_value_mux[5][9] , \read_value_mux[5][8] , \read_value_mux[5][7] , 
        \read_value_mux[5][6] , \read_value_mux[5][5] , \read_value_mux[5][4] , 
        \read_value_mux[5][3] , \read_value_mux[5][2] , \read_value_mux[5][1] , 
        \read_value_mux[5][0] , \read_value_mux[4][31] , 
        \read_value_mux[4][30] , \read_value_mux[4][29] , 
        \read_value_mux[4][28] , \read_value_mux[4][27] , 
        \read_value_mux[4][26] , \read_value_mux[4][25] , 
        \read_value_mux[4][24] , \read_value_mux[4][23] , 
        \read_value_mux[4][22] , \read_value_mux[4][21] , 
        \read_value_mux[4][20] , \read_value_mux[4][19] , 
        \read_value_mux[4][18] , \read_value_mux[4][17] , 
        \read_value_mux[4][16] , \read_value_mux[4][15] , 
        \read_value_mux[4][14] , \read_value_mux[4][13] , 
        \read_value_mux[4][12] , \read_value_mux[4][11] , 
        \read_value_mux[4][10] , \read_value_mux[4][9] , 
        \read_value_mux[4][8] , \read_value_mux[4][7] , \read_value_mux[4][6] , 
        \read_value_mux[4][5] , \read_value_mux[4][4] , \read_value_mux[4][3] , 
        \read_value_mux[4][2] , \read_value_mux[4][1] , \read_value_mux[4][0] , 
        \read_value_mux[3][31] , \read_value_mux[3][30] , 
        \read_value_mux[3][29] , \read_value_mux[3][28] , 
        \read_value_mux[3][27] , \read_value_mux[3][26] , 
        \read_value_mux[3][25] , \read_value_mux[3][24] , 
        \read_value_mux[3][23] , \read_value_mux[3][22] , 
        \read_value_mux[3][21] , \read_value_mux[3][20] , 
        \read_value_mux[3][19] , \read_value_mux[3][18] , 
        \read_value_mux[3][17] , \read_value_mux[3][16] , 
        \read_value_mux[3][15] , \read_value_mux[3][14] , 
        \read_value_mux[3][13] , \read_value_mux[3][12] , 
        \read_value_mux[3][11] , \read_value_mux[3][10] , 
        \read_value_mux[3][9] , \read_value_mux[3][8] , \read_value_mux[3][7] , 
        \read_value_mux[3][6] , \read_value_mux[3][5] , \read_value_mux[3][4] , 
        \read_value_mux[3][3] , \read_value_mux[3][2] , \read_value_mux[3][1] , 
        \read_value_mux[3][0] , \read_value_mux[2][31] , 
        \read_value_mux[2][30] , \read_value_mux[2][29] , 
        \read_value_mux[2][28] , \read_value_mux[2][27] , 
        \read_value_mux[2][26] , \read_value_mux[2][25] , 
        \read_value_mux[2][24] , \read_value_mux[2][23] , 
        \read_value_mux[2][22] , \read_value_mux[2][21] , 
        \read_value_mux[2][20] , \read_value_mux[2][19] , 
        \read_value_mux[2][18] , \read_value_mux[2][17] , 
        \read_value_mux[2][16] , \read_value_mux[2][15] , 
        \read_value_mux[2][14] , \read_value_mux[2][13] , 
        \read_value_mux[2][12] , \read_value_mux[2][11] , 
        \read_value_mux[2][10] , \read_value_mux[2][9] , 
        \read_value_mux[2][8] , \read_value_mux[2][7] , \read_value_mux[2][6] , 
        \read_value_mux[2][5] , \read_value_mux[2][4] , \read_value_mux[2][3] , 
        \read_value_mux[2][2] , \read_value_mux[2][1] , \read_value_mux[2][0] , 
        \read_value_mux[1][31] , \read_value_mux[1][30] , 
        \read_value_mux[1][29] , \read_value_mux[1][28] , 
        \read_value_mux[1][27] , \read_value_mux[1][26] , 
        \read_value_mux[1][25] , \read_value_mux[1][24] , 
        \read_value_mux[1][23] , \read_value_mux[1][22] , 
        \read_value_mux[1][21] , \read_value_mux[1][20] , 
        \read_value_mux[1][19] , \read_value_mux[1][18] , 
        \read_value_mux[1][17] , \read_value_mux[1][16] , 
        \read_value_mux[1][15] , \read_value_mux[1][14] , 
        \read_value_mux[1][13] , \read_value_mux[1][12] , 
        \read_value_mux[1][11] , \read_value_mux[1][10] , 
        \read_value_mux[1][9] , \read_value_mux[1][8] , \read_value_mux[1][7] , 
        \read_value_mux[1][6] , \read_value_mux[1][5] , \read_value_mux[1][4] , 
        \read_value_mux[1][3] , \read_value_mux[1][2] , \read_value_mux[1][1] , 
        \read_value_mux[1][0] , \read_value_mux[0][31] , 
        \read_value_mux[0][30] , \read_value_mux[0][29] , 
        \read_value_mux[0][28] , \read_value_mux[0][27] , 
        \read_value_mux[0][26] , \read_value_mux[0][25] , 
        \read_value_mux[0][24] , \read_value_mux[0][23] , 
        \read_value_mux[0][22] , \read_value_mux[0][21] , 
        \read_value_mux[0][20] , \read_value_mux[0][19] , 
        \read_value_mux[0][18] , \read_value_mux[0][17] , 
        \read_value_mux[0][16] , \read_value_mux[0][15] , 
        \read_value_mux[0][14] , \read_value_mux[0][13] , 
        \read_value_mux[0][12] , \read_value_mux[0][11] , 
        \read_value_mux[0][10] , \read_value_mux[0][9] , 
        \read_value_mux[0][8] , \read_value_mux[0][7] , \read_value_mux[0][6] , 
        \read_value_mux[0][5] , \read_value_mux[0][4] , \read_value_mux[0][3] , 
        \read_value_mux[0][2] , \read_value_mux[0][1] , \read_value_mux[0][0] }), .select_i(read_index), .data_o(read_value) );
  GTECH_OR2 C8 ( .A(N29), .B(read_results[0]), .Z(read_valid) );
  GTECH_OR2 C9 ( .A(N28), .B(read_results[1]), .Z(N29) );
  GTECH_OR2 C10 ( .A(N27), .B(read_results[2]), .Z(N28) );
  GTECH_OR2 C11 ( .A(N26), .B(read_results[3]), .Z(N27) );
  GTECH_OR2 C12 ( .A(N25), .B(read_results[4]), .Z(N26) );
  GTECH_OR2 C13 ( .A(N24), .B(read_results[5]), .Z(N25) );
  GTECH_OR2 C14 ( .A(N23), .B(read_results[6]), .Z(N24) );
  GTECH_OR2 C15 ( .A(N22), .B(read_results[7]), .Z(N23) );
  GTECH_OR2 C16 ( .A(N21), .B(read_results[8]), .Z(N22) );
  GTECH_OR2 C17 ( .A(N20), .B(read_results[9]), .Z(N21) );
  GTECH_OR2 C18 ( .A(N19), .B(read_results[10]), .Z(N20) );
  GTECH_OR2 C19 ( .A(N18), .B(read_results[11]), .Z(N19) );
  GTECH_OR2 C20 ( .A(N17), .B(read_results[12]), .Z(N18) );
  GTECH_OR2 C21 ( .A(N16), .B(read_results[13]), .Z(N17) );
  GTECH_OR2 C22 ( .A(N15), .B(read_results[14]), .Z(N16) );
  GTECH_OR2 C23 ( .A(N14), .B(read_results[15]), .Z(N15) );
  GTECH_OR2 C24 ( .A(N13), .B(read_results[16]), .Z(N14) );
  GTECH_OR2 C25 ( .A(N12), .B(read_results[17]), .Z(N13) );
  GTECH_OR2 C26 ( .A(N11), .B(read_results[18]), .Z(N12) );
  GTECH_OR2 C27 ( .A(N10), .B(read_results[19]), .Z(N11) );
  GTECH_OR2 C28 ( .A(N9), .B(read_results[20]), .Z(N10) );
  GTECH_OR2 C29 ( .A(N8), .B(read_results[21]), .Z(N9) );
  GTECH_OR2 C30 ( .A(N7), .B(read_results[22]), .Z(N8) );
  GTECH_OR2 C31 ( .A(N6), .B(read_results[23]), .Z(N7) );
  GTECH_OR2 C32 ( .A(N5), .B(read_results[24]), .Z(N6) );
  GTECH_OR2 C33 ( .A(N4), .B(read_results[25]), .Z(N5) );
  GTECH_OR2 C34 ( .A(N3), .B(read_results[26]), .Z(N4) );
  GTECH_OR2 C35 ( .A(N2), .B(read_results[27]), .Z(N3) );
  GTECH_OR2 C36 ( .A(N1), .B(read_results[28]), .Z(N2) );
  GTECH_OR2 C37 ( .A(N0), .B(read_results[29]), .Z(N1) );
  GTECH_OR2 C38 ( .A(read_results[31]), .B(read_results[30]), .Z(N0) );
  GTECH_OR2 C39 ( .A(N59), .B(search_results[0]), .Z(search_valid) );
  GTECH_OR2 C40 ( .A(N58), .B(search_results[1]), .Z(N59) );
  GTECH_OR2 C41 ( .A(N57), .B(search_results[2]), .Z(N58) );
  GTECH_OR2 C42 ( .A(N56), .B(search_results[3]), .Z(N57) );
  GTECH_OR2 C43 ( .A(N55), .B(search_results[4]), .Z(N56) );
  GTECH_OR2 C44 ( .A(N54), .B(search_results[5]), .Z(N55) );
  GTECH_OR2 C45 ( .A(N53), .B(search_results[6]), .Z(N54) );
  GTECH_OR2 C46 ( .A(N52), .B(search_results[7]), .Z(N53) );
  GTECH_OR2 C47 ( .A(N51), .B(search_results[8]), .Z(N52) );
  GTECH_OR2 C48 ( .A(N50), .B(search_results[9]), .Z(N51) );
  GTECH_OR2 C49 ( .A(N49), .B(search_results[10]), .Z(N50) );
  GTECH_OR2 C50 ( .A(N48), .B(search_results[11]), .Z(N49) );
  GTECH_OR2 C51 ( .A(N47), .B(search_results[12]), .Z(N48) );
  GTECH_OR2 C52 ( .A(N46), .B(search_results[13]), .Z(N47) );
  GTECH_OR2 C53 ( .A(N45), .B(search_results[14]), .Z(N46) );
  GTECH_OR2 C54 ( .A(N44), .B(search_results[15]), .Z(N45) );
  GTECH_OR2 C55 ( .A(N43), .B(search_results[16]), .Z(N44) );
  GTECH_OR2 C56 ( .A(N42), .B(search_results[17]), .Z(N43) );
  GTECH_OR2 C57 ( .A(N41), .B(search_results[18]), .Z(N42) );
  GTECH_OR2 C58 ( .A(N40), .B(search_results[19]), .Z(N41) );
  GTECH_OR2 C59 ( .A(N39), .B(search_results[20]), .Z(N40) );
  GTECH_OR2 C60 ( .A(N38), .B(search_results[21]), .Z(N39) );
  GTECH_OR2 C61 ( .A(N37), .B(search_results[22]), .Z(N38) );
  GTECH_OR2 C62 ( .A(N36), .B(search_results[23]), .Z(N37) );
  GTECH_OR2 C63 ( .A(N35), .B(search_results[24]), .Z(N36) );
  GTECH_OR2 C64 ( .A(N34), .B(search_results[25]), .Z(N35) );
  GTECH_OR2 C65 ( .A(N33), .B(search_results[26]), .Z(N34) );
  GTECH_OR2 C66 ( .A(N32), .B(search_results[27]), .Z(N33) );
  GTECH_OR2 C67 ( .A(N31), .B(search_results[28]), .Z(N32) );
  GTECH_OR2 C68 ( .A(N30), .B(search_results[29]), .Z(N31) );
  GTECH_OR2 C69 ( .A(search_results[31]), .B(search_results[30]), .Z(N30) );
endmodule

