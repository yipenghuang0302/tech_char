
module mux ( .data_i({\data_i[31][31] , \data_i[31][30] , \data_i[31][29] , 
        \data_i[31][28] , \data_i[31][27] , \data_i[31][26] , \data_i[31][25] , 
        \data_i[31][24] , \data_i[31][23] , \data_i[31][22] , \data_i[31][21] , 
        \data_i[31][20] , \data_i[31][19] , \data_i[31][18] , \data_i[31][17] , 
        \data_i[31][16] , \data_i[31][15] , \data_i[31][14] , \data_i[31][13] , 
        \data_i[31][12] , \data_i[31][11] , \data_i[31][10] , \data_i[31][9] , 
        \data_i[31][8] , \data_i[31][7] , \data_i[31][6] , \data_i[31][5] , 
        \data_i[31][4] , \data_i[31][3] , \data_i[31][2] , \data_i[31][1] , 
        \data_i[31][0] , \data_i[30][31] , \data_i[30][30] , \data_i[30][29] , 
        \data_i[30][28] , \data_i[30][27] , \data_i[30][26] , \data_i[30][25] , 
        \data_i[30][24] , \data_i[30][23] , \data_i[30][22] , \data_i[30][21] , 
        \data_i[30][20] , \data_i[30][19] , \data_i[30][18] , \data_i[30][17] , 
        \data_i[30][16] , \data_i[30][15] , \data_i[30][14] , \data_i[30][13] , 
        \data_i[30][12] , \data_i[30][11] , \data_i[30][10] , \data_i[30][9] , 
        \data_i[30][8] , \data_i[30][7] , \data_i[30][6] , \data_i[30][5] , 
        \data_i[30][4] , \data_i[30][3] , \data_i[30][2] , \data_i[30][1] , 
        \data_i[30][0] , \data_i[29][31] , \data_i[29][30] , \data_i[29][29] , 
        \data_i[29][28] , \data_i[29][27] , \data_i[29][26] , \data_i[29][25] , 
        \data_i[29][24] , \data_i[29][23] , \data_i[29][22] , \data_i[29][21] , 
        \data_i[29][20] , \data_i[29][19] , \data_i[29][18] , \data_i[29][17] , 
        \data_i[29][16] , \data_i[29][15] , \data_i[29][14] , \data_i[29][13] , 
        \data_i[29][12] , \data_i[29][11] , \data_i[29][10] , \data_i[29][9] , 
        \data_i[29][8] , \data_i[29][7] , \data_i[29][6] , \data_i[29][5] , 
        \data_i[29][4] , \data_i[29][3] , \data_i[29][2] , \data_i[29][1] , 
        \data_i[29][0] , \data_i[28][31] , \data_i[28][30] , \data_i[28][29] , 
        \data_i[28][28] , \data_i[28][27] , \data_i[28][26] , \data_i[28][25] , 
        \data_i[28][24] , \data_i[28][23] , \data_i[28][22] , \data_i[28][21] , 
        \data_i[28][20] , \data_i[28][19] , \data_i[28][18] , \data_i[28][17] , 
        \data_i[28][16] , \data_i[28][15] , \data_i[28][14] , \data_i[28][13] , 
        \data_i[28][12] , \data_i[28][11] , \data_i[28][10] , \data_i[28][9] , 
        \data_i[28][8] , \data_i[28][7] , \data_i[28][6] , \data_i[28][5] , 
        \data_i[28][4] , \data_i[28][3] , \data_i[28][2] , \data_i[28][1] , 
        \data_i[28][0] , \data_i[27][31] , \data_i[27][30] , \data_i[27][29] , 
        \data_i[27][28] , \data_i[27][27] , \data_i[27][26] , \data_i[27][25] , 
        \data_i[27][24] , \data_i[27][23] , \data_i[27][22] , \data_i[27][21] , 
        \data_i[27][20] , \data_i[27][19] , \data_i[27][18] , \data_i[27][17] , 
        \data_i[27][16] , \data_i[27][15] , \data_i[27][14] , \data_i[27][13] , 
        \data_i[27][12] , \data_i[27][11] , \data_i[27][10] , \data_i[27][9] , 
        \data_i[27][8] , \data_i[27][7] , \data_i[27][6] , \data_i[27][5] , 
        \data_i[27][4] , \data_i[27][3] , \data_i[27][2] , \data_i[27][1] , 
        \data_i[27][0] , \data_i[26][31] , \data_i[26][30] , \data_i[26][29] , 
        \data_i[26][28] , \data_i[26][27] , \data_i[26][26] , \data_i[26][25] , 
        \data_i[26][24] , \data_i[26][23] , \data_i[26][22] , \data_i[26][21] , 
        \data_i[26][20] , \data_i[26][19] , \data_i[26][18] , \data_i[26][17] , 
        \data_i[26][16] , \data_i[26][15] , \data_i[26][14] , \data_i[26][13] , 
        \data_i[26][12] , \data_i[26][11] , \data_i[26][10] , \data_i[26][9] , 
        \data_i[26][8] , \data_i[26][7] , \data_i[26][6] , \data_i[26][5] , 
        \data_i[26][4] , \data_i[26][3] , \data_i[26][2] , \data_i[26][1] , 
        \data_i[26][0] , \data_i[25][31] , \data_i[25][30] , \data_i[25][29] , 
        \data_i[25][28] , \data_i[25][27] , \data_i[25][26] , \data_i[25][25] , 
        \data_i[25][24] , \data_i[25][23] , \data_i[25][22] , \data_i[25][21] , 
        \data_i[25][20] , \data_i[25][19] , \data_i[25][18] , \data_i[25][17] , 
        \data_i[25][16] , \data_i[25][15] , \data_i[25][14] , \data_i[25][13] , 
        \data_i[25][12] , \data_i[25][11] , \data_i[25][10] , \data_i[25][9] , 
        \data_i[25][8] , \data_i[25][7] , \data_i[25][6] , \data_i[25][5] , 
        \data_i[25][4] , \data_i[25][3] , \data_i[25][2] , \data_i[25][1] , 
        \data_i[25][0] , \data_i[24][31] , \data_i[24][30] , \data_i[24][29] , 
        \data_i[24][28] , \data_i[24][27] , \data_i[24][26] , \data_i[24][25] , 
        \data_i[24][24] , \data_i[24][23] , \data_i[24][22] , \data_i[24][21] , 
        \data_i[24][20] , \data_i[24][19] , \data_i[24][18] , \data_i[24][17] , 
        \data_i[24][16] , \data_i[24][15] , \data_i[24][14] , \data_i[24][13] , 
        \data_i[24][12] , \data_i[24][11] , \data_i[24][10] , \data_i[24][9] , 
        \data_i[24][8] , \data_i[24][7] , \data_i[24][6] , \data_i[24][5] , 
        \data_i[24][4] , \data_i[24][3] , \data_i[24][2] , \data_i[24][1] , 
        \data_i[24][0] , \data_i[23][31] , \data_i[23][30] , \data_i[23][29] , 
        \data_i[23][28] , \data_i[23][27] , \data_i[23][26] , \data_i[23][25] , 
        \data_i[23][24] , \data_i[23][23] , \data_i[23][22] , \data_i[23][21] , 
        \data_i[23][20] , \data_i[23][19] , \data_i[23][18] , \data_i[23][17] , 
        \data_i[23][16] , \data_i[23][15] , \data_i[23][14] , \data_i[23][13] , 
        \data_i[23][12] , \data_i[23][11] , \data_i[23][10] , \data_i[23][9] , 
        \data_i[23][8] , \data_i[23][7] , \data_i[23][6] , \data_i[23][5] , 
        \data_i[23][4] , \data_i[23][3] , \data_i[23][2] , \data_i[23][1] , 
        \data_i[23][0] , \data_i[22][31] , \data_i[22][30] , \data_i[22][29] , 
        \data_i[22][28] , \data_i[22][27] , \data_i[22][26] , \data_i[22][25] , 
        \data_i[22][24] , \data_i[22][23] , \data_i[22][22] , \data_i[22][21] , 
        \data_i[22][20] , \data_i[22][19] , \data_i[22][18] , \data_i[22][17] , 
        \data_i[22][16] , \data_i[22][15] , \data_i[22][14] , \data_i[22][13] , 
        \data_i[22][12] , \data_i[22][11] , \data_i[22][10] , \data_i[22][9] , 
        \data_i[22][8] , \data_i[22][7] , \data_i[22][6] , \data_i[22][5] , 
        \data_i[22][4] , \data_i[22][3] , \data_i[22][2] , \data_i[22][1] , 
        \data_i[22][0] , \data_i[21][31] , \data_i[21][30] , \data_i[21][29] , 
        \data_i[21][28] , \data_i[21][27] , \data_i[21][26] , \data_i[21][25] , 
        \data_i[21][24] , \data_i[21][23] , \data_i[21][22] , \data_i[21][21] , 
        \data_i[21][20] , \data_i[21][19] , \data_i[21][18] , \data_i[21][17] , 
        \data_i[21][16] , \data_i[21][15] , \data_i[21][14] , \data_i[21][13] , 
        \data_i[21][12] , \data_i[21][11] , \data_i[21][10] , \data_i[21][9] , 
        \data_i[21][8] , \data_i[21][7] , \data_i[21][6] , \data_i[21][5] , 
        \data_i[21][4] , \data_i[21][3] , \data_i[21][2] , \data_i[21][1] , 
        \data_i[21][0] , \data_i[20][31] , \data_i[20][30] , \data_i[20][29] , 
        \data_i[20][28] , \data_i[20][27] , \data_i[20][26] , \data_i[20][25] , 
        \data_i[20][24] , \data_i[20][23] , \data_i[20][22] , \data_i[20][21] , 
        \data_i[20][20] , \data_i[20][19] , \data_i[20][18] , \data_i[20][17] , 
        \data_i[20][16] , \data_i[20][15] , \data_i[20][14] , \data_i[20][13] , 
        \data_i[20][12] , \data_i[20][11] , \data_i[20][10] , \data_i[20][9] , 
        \data_i[20][8] , \data_i[20][7] , \data_i[20][6] , \data_i[20][5] , 
        \data_i[20][4] , \data_i[20][3] , \data_i[20][2] , \data_i[20][1] , 
        \data_i[20][0] , \data_i[19][31] , \data_i[19][30] , \data_i[19][29] , 
        \data_i[19][28] , \data_i[19][27] , \data_i[19][26] , \data_i[19][25] , 
        \data_i[19][24] , \data_i[19][23] , \data_i[19][22] , \data_i[19][21] , 
        \data_i[19][20] , \data_i[19][19] , \data_i[19][18] , \data_i[19][17] , 
        \data_i[19][16] , \data_i[19][15] , \data_i[19][14] , \data_i[19][13] , 
        \data_i[19][12] , \data_i[19][11] , \data_i[19][10] , \data_i[19][9] , 
        \data_i[19][8] , \data_i[19][7] , \data_i[19][6] , \data_i[19][5] , 
        \data_i[19][4] , \data_i[19][3] , \data_i[19][2] , \data_i[19][1] , 
        \data_i[19][0] , \data_i[18][31] , \data_i[18][30] , \data_i[18][29] , 
        \data_i[18][28] , \data_i[18][27] , \data_i[18][26] , \data_i[18][25] , 
        \data_i[18][24] , \data_i[18][23] , \data_i[18][22] , \data_i[18][21] , 
        \data_i[18][20] , \data_i[18][19] , \data_i[18][18] , \data_i[18][17] , 
        \data_i[18][16] , \data_i[18][15] , \data_i[18][14] , \data_i[18][13] , 
        \data_i[18][12] , \data_i[18][11] , \data_i[18][10] , \data_i[18][9] , 
        \data_i[18][8] , \data_i[18][7] , \data_i[18][6] , \data_i[18][5] , 
        \data_i[18][4] , \data_i[18][3] , \data_i[18][2] , \data_i[18][1] , 
        \data_i[18][0] , \data_i[17][31] , \data_i[17][30] , \data_i[17][29] , 
        \data_i[17][28] , \data_i[17][27] , \data_i[17][26] , \data_i[17][25] , 
        \data_i[17][24] , \data_i[17][23] , \data_i[17][22] , \data_i[17][21] , 
        \data_i[17][20] , \data_i[17][19] , \data_i[17][18] , \data_i[17][17] , 
        \data_i[17][16] , \data_i[17][15] , \data_i[17][14] , \data_i[17][13] , 
        \data_i[17][12] , \data_i[17][11] , \data_i[17][10] , \data_i[17][9] , 
        \data_i[17][8] , \data_i[17][7] , \data_i[17][6] , \data_i[17][5] , 
        \data_i[17][4] , \data_i[17][3] , \data_i[17][2] , \data_i[17][1] , 
        \data_i[17][0] , \data_i[16][31] , \data_i[16][30] , \data_i[16][29] , 
        \data_i[16][28] , \data_i[16][27] , \data_i[16][26] , \data_i[16][25] , 
        \data_i[16][24] , \data_i[16][23] , \data_i[16][22] , \data_i[16][21] , 
        \data_i[16][20] , \data_i[16][19] , \data_i[16][18] , \data_i[16][17] , 
        \data_i[16][16] , \data_i[16][15] , \data_i[16][14] , \data_i[16][13] , 
        \data_i[16][12] , \data_i[16][11] , \data_i[16][10] , \data_i[16][9] , 
        \data_i[16][8] , \data_i[16][7] , \data_i[16][6] , \data_i[16][5] , 
        \data_i[16][4] , \data_i[16][3] , \data_i[16][2] , \data_i[16][1] , 
        \data_i[16][0] , \data_i[15][31] , \data_i[15][30] , \data_i[15][29] , 
        \data_i[15][28] , \data_i[15][27] , \data_i[15][26] , \data_i[15][25] , 
        \data_i[15][24] , \data_i[15][23] , \data_i[15][22] , \data_i[15][21] , 
        \data_i[15][20] , \data_i[15][19] , \data_i[15][18] , \data_i[15][17] , 
        \data_i[15][16] , \data_i[15][15] , \data_i[15][14] , \data_i[15][13] , 
        \data_i[15][12] , \data_i[15][11] , \data_i[15][10] , \data_i[15][9] , 
        \data_i[15][8] , \data_i[15][7] , \data_i[15][6] , \data_i[15][5] , 
        \data_i[15][4] , \data_i[15][3] , \data_i[15][2] , \data_i[15][1] , 
        \data_i[15][0] , \data_i[14][31] , \data_i[14][30] , \data_i[14][29] , 
        \data_i[14][28] , \data_i[14][27] , \data_i[14][26] , \data_i[14][25] , 
        \data_i[14][24] , \data_i[14][23] , \data_i[14][22] , \data_i[14][21] , 
        \data_i[14][20] , \data_i[14][19] , \data_i[14][18] , \data_i[14][17] , 
        \data_i[14][16] , \data_i[14][15] , \data_i[14][14] , \data_i[14][13] , 
        \data_i[14][12] , \data_i[14][11] , \data_i[14][10] , \data_i[14][9] , 
        \data_i[14][8] , \data_i[14][7] , \data_i[14][6] , \data_i[14][5] , 
        \data_i[14][4] , \data_i[14][3] , \data_i[14][2] , \data_i[14][1] , 
        \data_i[14][0] , \data_i[13][31] , \data_i[13][30] , \data_i[13][29] , 
        \data_i[13][28] , \data_i[13][27] , \data_i[13][26] , \data_i[13][25] , 
        \data_i[13][24] , \data_i[13][23] , \data_i[13][22] , \data_i[13][21] , 
        \data_i[13][20] , \data_i[13][19] , \data_i[13][18] , \data_i[13][17] , 
        \data_i[13][16] , \data_i[13][15] , \data_i[13][14] , \data_i[13][13] , 
        \data_i[13][12] , \data_i[13][11] , \data_i[13][10] , \data_i[13][9] , 
        \data_i[13][8] , \data_i[13][7] , \data_i[13][6] , \data_i[13][5] , 
        \data_i[13][4] , \data_i[13][3] , \data_i[13][2] , \data_i[13][1] , 
        \data_i[13][0] , \data_i[12][31] , \data_i[12][30] , \data_i[12][29] , 
        \data_i[12][28] , \data_i[12][27] , \data_i[12][26] , \data_i[12][25] , 
        \data_i[12][24] , \data_i[12][23] , \data_i[12][22] , \data_i[12][21] , 
        \data_i[12][20] , \data_i[12][19] , \data_i[12][18] , \data_i[12][17] , 
        \data_i[12][16] , \data_i[12][15] , \data_i[12][14] , \data_i[12][13] , 
        \data_i[12][12] , \data_i[12][11] , \data_i[12][10] , \data_i[12][9] , 
        \data_i[12][8] , \data_i[12][7] , \data_i[12][6] , \data_i[12][5] , 
        \data_i[12][4] , \data_i[12][3] , \data_i[12][2] , \data_i[12][1] , 
        \data_i[12][0] , \data_i[11][31] , \data_i[11][30] , \data_i[11][29] , 
        \data_i[11][28] , \data_i[11][27] , \data_i[11][26] , \data_i[11][25] , 
        \data_i[11][24] , \data_i[11][23] , \data_i[11][22] , \data_i[11][21] , 
        \data_i[11][20] , \data_i[11][19] , \data_i[11][18] , \data_i[11][17] , 
        \data_i[11][16] , \data_i[11][15] , \data_i[11][14] , \data_i[11][13] , 
        \data_i[11][12] , \data_i[11][11] , \data_i[11][10] , \data_i[11][9] , 
        \data_i[11][8] , \data_i[11][7] , \data_i[11][6] , \data_i[11][5] , 
        \data_i[11][4] , \data_i[11][3] , \data_i[11][2] , \data_i[11][1] , 
        \data_i[11][0] , \data_i[10][31] , \data_i[10][30] , \data_i[10][29] , 
        \data_i[10][28] , \data_i[10][27] , \data_i[10][26] , \data_i[10][25] , 
        \data_i[10][24] , \data_i[10][23] , \data_i[10][22] , \data_i[10][21] , 
        \data_i[10][20] , \data_i[10][19] , \data_i[10][18] , \data_i[10][17] , 
        \data_i[10][16] , \data_i[10][15] , \data_i[10][14] , \data_i[10][13] , 
        \data_i[10][12] , \data_i[10][11] , \data_i[10][10] , \data_i[10][9] , 
        \data_i[10][8] , \data_i[10][7] , \data_i[10][6] , \data_i[10][5] , 
        \data_i[10][4] , \data_i[10][3] , \data_i[10][2] , \data_i[10][1] , 
        \data_i[10][0] , \data_i[9][31] , \data_i[9][30] , \data_i[9][29] , 
        \data_i[9][28] , \data_i[9][27] , \data_i[9][26] , \data_i[9][25] , 
        \data_i[9][24] , \data_i[9][23] , \data_i[9][22] , \data_i[9][21] , 
        \data_i[9][20] , \data_i[9][19] , \data_i[9][18] , \data_i[9][17] , 
        \data_i[9][16] , \data_i[9][15] , \data_i[9][14] , \data_i[9][13] , 
        \data_i[9][12] , \data_i[9][11] , \data_i[9][10] , \data_i[9][9] , 
        \data_i[9][8] , \data_i[9][7] , \data_i[9][6] , \data_i[9][5] , 
        \data_i[9][4] , \data_i[9][3] , \data_i[9][2] , \data_i[9][1] , 
        \data_i[9][0] , \data_i[8][31] , \data_i[8][30] , \data_i[8][29] , 
        \data_i[8][28] , \data_i[8][27] , \data_i[8][26] , \data_i[8][25] , 
        \data_i[8][24] , \data_i[8][23] , \data_i[8][22] , \data_i[8][21] , 
        \data_i[8][20] , \data_i[8][19] , \data_i[8][18] , \data_i[8][17] , 
        \data_i[8][16] , \data_i[8][15] , \data_i[8][14] , \data_i[8][13] , 
        \data_i[8][12] , \data_i[8][11] , \data_i[8][10] , \data_i[8][9] , 
        \data_i[8][8] , \data_i[8][7] , \data_i[8][6] , \data_i[8][5] , 
        \data_i[8][4] , \data_i[8][3] , \data_i[8][2] , \data_i[8][1] , 
        \data_i[8][0] , \data_i[7][31] , \data_i[7][30] , \data_i[7][29] , 
        \data_i[7][28] , \data_i[7][27] , \data_i[7][26] , \data_i[7][25] , 
        \data_i[7][24] , \data_i[7][23] , \data_i[7][22] , \data_i[7][21] , 
        \data_i[7][20] , \data_i[7][19] , \data_i[7][18] , \data_i[7][17] , 
        \data_i[7][16] , \data_i[7][15] , \data_i[7][14] , \data_i[7][13] , 
        \data_i[7][12] , \data_i[7][11] , \data_i[7][10] , \data_i[7][9] , 
        \data_i[7][8] , \data_i[7][7] , \data_i[7][6] , \data_i[7][5] , 
        \data_i[7][4] , \data_i[7][3] , \data_i[7][2] , \data_i[7][1] , 
        \data_i[7][0] , \data_i[6][31] , \data_i[6][30] , \data_i[6][29] , 
        \data_i[6][28] , \data_i[6][27] , \data_i[6][26] , \data_i[6][25] , 
        \data_i[6][24] , \data_i[6][23] , \data_i[6][22] , \data_i[6][21] , 
        \data_i[6][20] , \data_i[6][19] , \data_i[6][18] , \data_i[6][17] , 
        \data_i[6][16] , \data_i[6][15] , \data_i[6][14] , \data_i[6][13] , 
        \data_i[6][12] , \data_i[6][11] , \data_i[6][10] , \data_i[6][9] , 
        \data_i[6][8] , \data_i[6][7] , \data_i[6][6] , \data_i[6][5] , 
        \data_i[6][4] , \data_i[6][3] , \data_i[6][2] , \data_i[6][1] , 
        \data_i[6][0] , \data_i[5][31] , \data_i[5][30] , \data_i[5][29] , 
        \data_i[5][28] , \data_i[5][27] , \data_i[5][26] , \data_i[5][25] , 
        \data_i[5][24] , \data_i[5][23] , \data_i[5][22] , \data_i[5][21] , 
        \data_i[5][20] , \data_i[5][19] , \data_i[5][18] , \data_i[5][17] , 
        \data_i[5][16] , \data_i[5][15] , \data_i[5][14] , \data_i[5][13] , 
        \data_i[5][12] , \data_i[5][11] , \data_i[5][10] , \data_i[5][9] , 
        \data_i[5][8] , \data_i[5][7] , \data_i[5][6] , \data_i[5][5] , 
        \data_i[5][4] , \data_i[5][3] , \data_i[5][2] , \data_i[5][1] , 
        \data_i[5][0] , \data_i[4][31] , \data_i[4][30] , \data_i[4][29] , 
        \data_i[4][28] , \data_i[4][27] , \data_i[4][26] , \data_i[4][25] , 
        \data_i[4][24] , \data_i[4][23] , \data_i[4][22] , \data_i[4][21] , 
        \data_i[4][20] , \data_i[4][19] , \data_i[4][18] , \data_i[4][17] , 
        \data_i[4][16] , \data_i[4][15] , \data_i[4][14] , \data_i[4][13] , 
        \data_i[4][12] , \data_i[4][11] , \data_i[4][10] , \data_i[4][9] , 
        \data_i[4][8] , \data_i[4][7] , \data_i[4][6] , \data_i[4][5] , 
        \data_i[4][4] , \data_i[4][3] , \data_i[4][2] , \data_i[4][1] , 
        \data_i[4][0] , \data_i[3][31] , \data_i[3][30] , \data_i[3][29] , 
        \data_i[3][28] , \data_i[3][27] , \data_i[3][26] , \data_i[3][25] , 
        \data_i[3][24] , \data_i[3][23] , \data_i[3][22] , \data_i[3][21] , 
        \data_i[3][20] , \data_i[3][19] , \data_i[3][18] , \data_i[3][17] , 
        \data_i[3][16] , \data_i[3][15] , \data_i[3][14] , \data_i[3][13] , 
        \data_i[3][12] , \data_i[3][11] , \data_i[3][10] , \data_i[3][9] , 
        \data_i[3][8] , \data_i[3][7] , \data_i[3][6] , \data_i[3][5] , 
        \data_i[3][4] , \data_i[3][3] , \data_i[3][2] , \data_i[3][1] , 
        \data_i[3][0] , \data_i[2][31] , \data_i[2][30] , \data_i[2][29] , 
        \data_i[2][28] , \data_i[2][27] , \data_i[2][26] , \data_i[2][25] , 
        \data_i[2][24] , \data_i[2][23] , \data_i[2][22] , \data_i[2][21] , 
        \data_i[2][20] , \data_i[2][19] , \data_i[2][18] , \data_i[2][17] , 
        \data_i[2][16] , \data_i[2][15] , \data_i[2][14] , \data_i[2][13] , 
        \data_i[2][12] , \data_i[2][11] , \data_i[2][10] , \data_i[2][9] , 
        \data_i[2][8] , \data_i[2][7] , \data_i[2][6] , \data_i[2][5] , 
        \data_i[2][4] , \data_i[2][3] , \data_i[2][2] , \data_i[2][1] , 
        \data_i[2][0] , \data_i[1][31] , \data_i[1][30] , \data_i[1][29] , 
        \data_i[1][28] , \data_i[1][27] , \data_i[1][26] , \data_i[1][25] , 
        \data_i[1][24] , \data_i[1][23] , \data_i[1][22] , \data_i[1][21] , 
        \data_i[1][20] , \data_i[1][19] , \data_i[1][18] , \data_i[1][17] , 
        \data_i[1][16] , \data_i[1][15] , \data_i[1][14] , \data_i[1][13] , 
        \data_i[1][12] , \data_i[1][11] , \data_i[1][10] , \data_i[1][9] , 
        \data_i[1][8] , \data_i[1][7] , \data_i[1][6] , \data_i[1][5] , 
        \data_i[1][4] , \data_i[1][3] , \data_i[1][2] , \data_i[1][1] , 
        \data_i[1][0] , \data_i[0][31] , \data_i[0][30] , \data_i[0][29] , 
        \data_i[0][28] , \data_i[0][27] , \data_i[0][26] , \data_i[0][25] , 
        \data_i[0][24] , \data_i[0][23] , \data_i[0][22] , \data_i[0][21] , 
        \data_i[0][20] , \data_i[0][19] , \data_i[0][18] , \data_i[0][17] , 
        \data_i[0][16] , \data_i[0][15] , \data_i[0][14] , \data_i[0][13] , 
        \data_i[0][12] , \data_i[0][11] , \data_i[0][10] , \data_i[0][9] , 
        \data_i[0][8] , \data_i[0][7] , \data_i[0][6] , \data_i[0][5] , 
        \data_i[0][4] , \data_i[0][3] , \data_i[0][2] , \data_i[0][1] , 
        \data_i[0][0] }), select_i, data_o );
  input [4:0] select_i;
  output [31:0] data_o;
  input \data_i[31][31] , \data_i[31][30] , \data_i[31][29] , \data_i[31][28] ,
         \data_i[31][27] , \data_i[31][26] , \data_i[31][25] ,
         \data_i[31][24] , \data_i[31][23] , \data_i[31][22] ,
         \data_i[31][21] , \data_i[31][20] , \data_i[31][19] ,
         \data_i[31][18] , \data_i[31][17] , \data_i[31][16] ,
         \data_i[31][15] , \data_i[31][14] , \data_i[31][13] ,
         \data_i[31][12] , \data_i[31][11] , \data_i[31][10] , \data_i[31][9] ,
         \data_i[31][8] , \data_i[31][7] , \data_i[31][6] , \data_i[31][5] ,
         \data_i[31][4] , \data_i[31][3] , \data_i[31][2] , \data_i[31][1] ,
         \data_i[31][0] , \data_i[30][31] , \data_i[30][30] , \data_i[30][29] ,
         \data_i[30][28] , \data_i[30][27] , \data_i[30][26] ,
         \data_i[30][25] , \data_i[30][24] , \data_i[30][23] ,
         \data_i[30][22] , \data_i[30][21] , \data_i[30][20] ,
         \data_i[30][19] , \data_i[30][18] , \data_i[30][17] ,
         \data_i[30][16] , \data_i[30][15] , \data_i[30][14] ,
         \data_i[30][13] , \data_i[30][12] , \data_i[30][11] ,
         \data_i[30][10] , \data_i[30][9] , \data_i[30][8] , \data_i[30][7] ,
         \data_i[30][6] , \data_i[30][5] , \data_i[30][4] , \data_i[30][3] ,
         \data_i[30][2] , \data_i[30][1] , \data_i[30][0] , \data_i[29][31] ,
         \data_i[29][30] , \data_i[29][29] , \data_i[29][28] ,
         \data_i[29][27] , \data_i[29][26] , \data_i[29][25] ,
         \data_i[29][24] , \data_i[29][23] , \data_i[29][22] ,
         \data_i[29][21] , \data_i[29][20] , \data_i[29][19] ,
         \data_i[29][18] , \data_i[29][17] , \data_i[29][16] ,
         \data_i[29][15] , \data_i[29][14] , \data_i[29][13] ,
         \data_i[29][12] , \data_i[29][11] , \data_i[29][10] , \data_i[29][9] ,
         \data_i[29][8] , \data_i[29][7] , \data_i[29][6] , \data_i[29][5] ,
         \data_i[29][4] , \data_i[29][3] , \data_i[29][2] , \data_i[29][1] ,
         \data_i[29][0] , \data_i[28][31] , \data_i[28][30] , \data_i[28][29] ,
         \data_i[28][28] , \data_i[28][27] , \data_i[28][26] ,
         \data_i[28][25] , \data_i[28][24] , \data_i[28][23] ,
         \data_i[28][22] , \data_i[28][21] , \data_i[28][20] ,
         \data_i[28][19] , \data_i[28][18] , \data_i[28][17] ,
         \data_i[28][16] , \data_i[28][15] , \data_i[28][14] ,
         \data_i[28][13] , \data_i[28][12] , \data_i[28][11] ,
         \data_i[28][10] , \data_i[28][9] , \data_i[28][8] , \data_i[28][7] ,
         \data_i[28][6] , \data_i[28][5] , \data_i[28][4] , \data_i[28][3] ,
         \data_i[28][2] , \data_i[28][1] , \data_i[28][0] , \data_i[27][31] ,
         \data_i[27][30] , \data_i[27][29] , \data_i[27][28] ,
         \data_i[27][27] , \data_i[27][26] , \data_i[27][25] ,
         \data_i[27][24] , \data_i[27][23] , \data_i[27][22] ,
         \data_i[27][21] , \data_i[27][20] , \data_i[27][19] ,
         \data_i[27][18] , \data_i[27][17] , \data_i[27][16] ,
         \data_i[27][15] , \data_i[27][14] , \data_i[27][13] ,
         \data_i[27][12] , \data_i[27][11] , \data_i[27][10] , \data_i[27][9] ,
         \data_i[27][8] , \data_i[27][7] , \data_i[27][6] , \data_i[27][5] ,
         \data_i[27][4] , \data_i[27][3] , \data_i[27][2] , \data_i[27][1] ,
         \data_i[27][0] , \data_i[26][31] , \data_i[26][30] , \data_i[26][29] ,
         \data_i[26][28] , \data_i[26][27] , \data_i[26][26] ,
         \data_i[26][25] , \data_i[26][24] , \data_i[26][23] ,
         \data_i[26][22] , \data_i[26][21] , \data_i[26][20] ,
         \data_i[26][19] , \data_i[26][18] , \data_i[26][17] ,
         \data_i[26][16] , \data_i[26][15] , \data_i[26][14] ,
         \data_i[26][13] , \data_i[26][12] , \data_i[26][11] ,
         \data_i[26][10] , \data_i[26][9] , \data_i[26][8] , \data_i[26][7] ,
         \data_i[26][6] , \data_i[26][5] , \data_i[26][4] , \data_i[26][3] ,
         \data_i[26][2] , \data_i[26][1] , \data_i[26][0] , \data_i[25][31] ,
         \data_i[25][30] , \data_i[25][29] , \data_i[25][28] ,
         \data_i[25][27] , \data_i[25][26] , \data_i[25][25] ,
         \data_i[25][24] , \data_i[25][23] , \data_i[25][22] ,
         \data_i[25][21] , \data_i[25][20] , \data_i[25][19] ,
         \data_i[25][18] , \data_i[25][17] , \data_i[25][16] ,
         \data_i[25][15] , \data_i[25][14] , \data_i[25][13] ,
         \data_i[25][12] , \data_i[25][11] , \data_i[25][10] , \data_i[25][9] ,
         \data_i[25][8] , \data_i[25][7] , \data_i[25][6] , \data_i[25][5] ,
         \data_i[25][4] , \data_i[25][3] , \data_i[25][2] , \data_i[25][1] ,
         \data_i[25][0] , \data_i[24][31] , \data_i[24][30] , \data_i[24][29] ,
         \data_i[24][28] , \data_i[24][27] , \data_i[24][26] ,
         \data_i[24][25] , \data_i[24][24] , \data_i[24][23] ,
         \data_i[24][22] , \data_i[24][21] , \data_i[24][20] ,
         \data_i[24][19] , \data_i[24][18] , \data_i[24][17] ,
         \data_i[24][16] , \data_i[24][15] , \data_i[24][14] ,
         \data_i[24][13] , \data_i[24][12] , \data_i[24][11] ,
         \data_i[24][10] , \data_i[24][9] , \data_i[24][8] , \data_i[24][7] ,
         \data_i[24][6] , \data_i[24][5] , \data_i[24][4] , \data_i[24][3] ,
         \data_i[24][2] , \data_i[24][1] , \data_i[24][0] , \data_i[23][31] ,
         \data_i[23][30] , \data_i[23][29] , \data_i[23][28] ,
         \data_i[23][27] , \data_i[23][26] , \data_i[23][25] ,
         \data_i[23][24] , \data_i[23][23] , \data_i[23][22] ,
         \data_i[23][21] , \data_i[23][20] , \data_i[23][19] ,
         \data_i[23][18] , \data_i[23][17] , \data_i[23][16] ,
         \data_i[23][15] , \data_i[23][14] , \data_i[23][13] ,
         \data_i[23][12] , \data_i[23][11] , \data_i[23][10] , \data_i[23][9] ,
         \data_i[23][8] , \data_i[23][7] , \data_i[23][6] , \data_i[23][5] ,
         \data_i[23][4] , \data_i[23][3] , \data_i[23][2] , \data_i[23][1] ,
         \data_i[23][0] , \data_i[22][31] , \data_i[22][30] , \data_i[22][29] ,
         \data_i[22][28] , \data_i[22][27] , \data_i[22][26] ,
         \data_i[22][25] , \data_i[22][24] , \data_i[22][23] ,
         \data_i[22][22] , \data_i[22][21] , \data_i[22][20] ,
         \data_i[22][19] , \data_i[22][18] , \data_i[22][17] ,
         \data_i[22][16] , \data_i[22][15] , \data_i[22][14] ,
         \data_i[22][13] , \data_i[22][12] , \data_i[22][11] ,
         \data_i[22][10] , \data_i[22][9] , \data_i[22][8] , \data_i[22][7] ,
         \data_i[22][6] , \data_i[22][5] , \data_i[22][4] , \data_i[22][3] ,
         \data_i[22][2] , \data_i[22][1] , \data_i[22][0] , \data_i[21][31] ,
         \data_i[21][30] , \data_i[21][29] , \data_i[21][28] ,
         \data_i[21][27] , \data_i[21][26] , \data_i[21][25] ,
         \data_i[21][24] , \data_i[21][23] , \data_i[21][22] ,
         \data_i[21][21] , \data_i[21][20] , \data_i[21][19] ,
         \data_i[21][18] , \data_i[21][17] , \data_i[21][16] ,
         \data_i[21][15] , \data_i[21][14] , \data_i[21][13] ,
         \data_i[21][12] , \data_i[21][11] , \data_i[21][10] , \data_i[21][9] ,
         \data_i[21][8] , \data_i[21][7] , \data_i[21][6] , \data_i[21][5] ,
         \data_i[21][4] , \data_i[21][3] , \data_i[21][2] , \data_i[21][1] ,
         \data_i[21][0] , \data_i[20][31] , \data_i[20][30] , \data_i[20][29] ,
         \data_i[20][28] , \data_i[20][27] , \data_i[20][26] ,
         \data_i[20][25] , \data_i[20][24] , \data_i[20][23] ,
         \data_i[20][22] , \data_i[20][21] , \data_i[20][20] ,
         \data_i[20][19] , \data_i[20][18] , \data_i[20][17] ,
         \data_i[20][16] , \data_i[20][15] , \data_i[20][14] ,
         \data_i[20][13] , \data_i[20][12] , \data_i[20][11] ,
         \data_i[20][10] , \data_i[20][9] , \data_i[20][8] , \data_i[20][7] ,
         \data_i[20][6] , \data_i[20][5] , \data_i[20][4] , \data_i[20][3] ,
         \data_i[20][2] , \data_i[20][1] , \data_i[20][0] , \data_i[19][31] ,
         \data_i[19][30] , \data_i[19][29] , \data_i[19][28] ,
         \data_i[19][27] , \data_i[19][26] , \data_i[19][25] ,
         \data_i[19][24] , \data_i[19][23] , \data_i[19][22] ,
         \data_i[19][21] , \data_i[19][20] , \data_i[19][19] ,
         \data_i[19][18] , \data_i[19][17] , \data_i[19][16] ,
         \data_i[19][15] , \data_i[19][14] , \data_i[19][13] ,
         \data_i[19][12] , \data_i[19][11] , \data_i[19][10] , \data_i[19][9] ,
         \data_i[19][8] , \data_i[19][7] , \data_i[19][6] , \data_i[19][5] ,
         \data_i[19][4] , \data_i[19][3] , \data_i[19][2] , \data_i[19][1] ,
         \data_i[19][0] , \data_i[18][31] , \data_i[18][30] , \data_i[18][29] ,
         \data_i[18][28] , \data_i[18][27] , \data_i[18][26] ,
         \data_i[18][25] , \data_i[18][24] , \data_i[18][23] ,
         \data_i[18][22] , \data_i[18][21] , \data_i[18][20] ,
         \data_i[18][19] , \data_i[18][18] , \data_i[18][17] ,
         \data_i[18][16] , \data_i[18][15] , \data_i[18][14] ,
         \data_i[18][13] , \data_i[18][12] , \data_i[18][11] ,
         \data_i[18][10] , \data_i[18][9] , \data_i[18][8] , \data_i[18][7] ,
         \data_i[18][6] , \data_i[18][5] , \data_i[18][4] , \data_i[18][3] ,
         \data_i[18][2] , \data_i[18][1] , \data_i[18][0] , \data_i[17][31] ,
         \data_i[17][30] , \data_i[17][29] , \data_i[17][28] ,
         \data_i[17][27] , \data_i[17][26] , \data_i[17][25] ,
         \data_i[17][24] , \data_i[17][23] , \data_i[17][22] ,
         \data_i[17][21] , \data_i[17][20] , \data_i[17][19] ,
         \data_i[17][18] , \data_i[17][17] , \data_i[17][16] ,
         \data_i[17][15] , \data_i[17][14] , \data_i[17][13] ,
         \data_i[17][12] , \data_i[17][11] , \data_i[17][10] , \data_i[17][9] ,
         \data_i[17][8] , \data_i[17][7] , \data_i[17][6] , \data_i[17][5] ,
         \data_i[17][4] , \data_i[17][3] , \data_i[17][2] , \data_i[17][1] ,
         \data_i[17][0] , \data_i[16][31] , \data_i[16][30] , \data_i[16][29] ,
         \data_i[16][28] , \data_i[16][27] , \data_i[16][26] ,
         \data_i[16][25] , \data_i[16][24] , \data_i[16][23] ,
         \data_i[16][22] , \data_i[16][21] , \data_i[16][20] ,
         \data_i[16][19] , \data_i[16][18] , \data_i[16][17] ,
         \data_i[16][16] , \data_i[16][15] , \data_i[16][14] ,
         \data_i[16][13] , \data_i[16][12] , \data_i[16][11] ,
         \data_i[16][10] , \data_i[16][9] , \data_i[16][8] , \data_i[16][7] ,
         \data_i[16][6] , \data_i[16][5] , \data_i[16][4] , \data_i[16][3] ,
         \data_i[16][2] , \data_i[16][1] , \data_i[16][0] , \data_i[15][31] ,
         \data_i[15][30] , \data_i[15][29] , \data_i[15][28] ,
         \data_i[15][27] , \data_i[15][26] , \data_i[15][25] ,
         \data_i[15][24] , \data_i[15][23] , \data_i[15][22] ,
         \data_i[15][21] , \data_i[15][20] , \data_i[15][19] ,
         \data_i[15][18] , \data_i[15][17] , \data_i[15][16] ,
         \data_i[15][15] , \data_i[15][14] , \data_i[15][13] ,
         \data_i[15][12] , \data_i[15][11] , \data_i[15][10] , \data_i[15][9] ,
         \data_i[15][8] , \data_i[15][7] , \data_i[15][6] , \data_i[15][5] ,
         \data_i[15][4] , \data_i[15][3] , \data_i[15][2] , \data_i[15][1] ,
         \data_i[15][0] , \data_i[14][31] , \data_i[14][30] , \data_i[14][29] ,
         \data_i[14][28] , \data_i[14][27] , \data_i[14][26] ,
         \data_i[14][25] , \data_i[14][24] , \data_i[14][23] ,
         \data_i[14][22] , \data_i[14][21] , \data_i[14][20] ,
         \data_i[14][19] , \data_i[14][18] , \data_i[14][17] ,
         \data_i[14][16] , \data_i[14][15] , \data_i[14][14] ,
         \data_i[14][13] , \data_i[14][12] , \data_i[14][11] ,
         \data_i[14][10] , \data_i[14][9] , \data_i[14][8] , \data_i[14][7] ,
         \data_i[14][6] , \data_i[14][5] , \data_i[14][4] , \data_i[14][3] ,
         \data_i[14][2] , \data_i[14][1] , \data_i[14][0] , \data_i[13][31] ,
         \data_i[13][30] , \data_i[13][29] , \data_i[13][28] ,
         \data_i[13][27] , \data_i[13][26] , \data_i[13][25] ,
         \data_i[13][24] , \data_i[13][23] , \data_i[13][22] ,
         \data_i[13][21] , \data_i[13][20] , \data_i[13][19] ,
         \data_i[13][18] , \data_i[13][17] , \data_i[13][16] ,
         \data_i[13][15] , \data_i[13][14] , \data_i[13][13] ,
         \data_i[13][12] , \data_i[13][11] , \data_i[13][10] , \data_i[13][9] ,
         \data_i[13][8] , \data_i[13][7] , \data_i[13][6] , \data_i[13][5] ,
         \data_i[13][4] , \data_i[13][3] , \data_i[13][2] , \data_i[13][1] ,
         \data_i[13][0] , \data_i[12][31] , \data_i[12][30] , \data_i[12][29] ,
         \data_i[12][28] , \data_i[12][27] , \data_i[12][26] ,
         \data_i[12][25] , \data_i[12][24] , \data_i[12][23] ,
         \data_i[12][22] , \data_i[12][21] , \data_i[12][20] ,
         \data_i[12][19] , \data_i[12][18] , \data_i[12][17] ,
         \data_i[12][16] , \data_i[12][15] , \data_i[12][14] ,
         \data_i[12][13] , \data_i[12][12] , \data_i[12][11] ,
         \data_i[12][10] , \data_i[12][9] , \data_i[12][8] , \data_i[12][7] ,
         \data_i[12][6] , \data_i[12][5] , \data_i[12][4] , \data_i[12][3] ,
         \data_i[12][2] , \data_i[12][1] , \data_i[12][0] , \data_i[11][31] ,
         \data_i[11][30] , \data_i[11][29] , \data_i[11][28] ,
         \data_i[11][27] , \data_i[11][26] , \data_i[11][25] ,
         \data_i[11][24] , \data_i[11][23] , \data_i[11][22] ,
         \data_i[11][21] , \data_i[11][20] , \data_i[11][19] ,
         \data_i[11][18] , \data_i[11][17] , \data_i[11][16] ,
         \data_i[11][15] , \data_i[11][14] , \data_i[11][13] ,
         \data_i[11][12] , \data_i[11][11] , \data_i[11][10] , \data_i[11][9] ,
         \data_i[11][8] , \data_i[11][7] , \data_i[11][6] , \data_i[11][5] ,
         \data_i[11][4] , \data_i[11][3] , \data_i[11][2] , \data_i[11][1] ,
         \data_i[11][0] , \data_i[10][31] , \data_i[10][30] , \data_i[10][29] ,
         \data_i[10][28] , \data_i[10][27] , \data_i[10][26] ,
         \data_i[10][25] , \data_i[10][24] , \data_i[10][23] ,
         \data_i[10][22] , \data_i[10][21] , \data_i[10][20] ,
         \data_i[10][19] , \data_i[10][18] , \data_i[10][17] ,
         \data_i[10][16] , \data_i[10][15] , \data_i[10][14] ,
         \data_i[10][13] , \data_i[10][12] , \data_i[10][11] ,
         \data_i[10][10] , \data_i[10][9] , \data_i[10][8] , \data_i[10][7] ,
         \data_i[10][6] , \data_i[10][5] , \data_i[10][4] , \data_i[10][3] ,
         \data_i[10][2] , \data_i[10][1] , \data_i[10][0] , \data_i[9][31] ,
         \data_i[9][30] , \data_i[9][29] , \data_i[9][28] , \data_i[9][27] ,
         \data_i[9][26] , \data_i[9][25] , \data_i[9][24] , \data_i[9][23] ,
         \data_i[9][22] , \data_i[9][21] , \data_i[9][20] , \data_i[9][19] ,
         \data_i[9][18] , \data_i[9][17] , \data_i[9][16] , \data_i[9][15] ,
         \data_i[9][14] , \data_i[9][13] , \data_i[9][12] , \data_i[9][11] ,
         \data_i[9][10] , \data_i[9][9] , \data_i[9][8] , \data_i[9][7] ,
         \data_i[9][6] , \data_i[9][5] , \data_i[9][4] , \data_i[9][3] ,
         \data_i[9][2] , \data_i[9][1] , \data_i[9][0] , \data_i[8][31] ,
         \data_i[8][30] , \data_i[8][29] , \data_i[8][28] , \data_i[8][27] ,
         \data_i[8][26] , \data_i[8][25] , \data_i[8][24] , \data_i[8][23] ,
         \data_i[8][22] , \data_i[8][21] , \data_i[8][20] , \data_i[8][19] ,
         \data_i[8][18] , \data_i[8][17] , \data_i[8][16] , \data_i[8][15] ,
         \data_i[8][14] , \data_i[8][13] , \data_i[8][12] , \data_i[8][11] ,
         \data_i[8][10] , \data_i[8][9] , \data_i[8][8] , \data_i[8][7] ,
         \data_i[8][6] , \data_i[8][5] , \data_i[8][4] , \data_i[8][3] ,
         \data_i[8][2] , \data_i[8][1] , \data_i[8][0] , \data_i[7][31] ,
         \data_i[7][30] , \data_i[7][29] , \data_i[7][28] , \data_i[7][27] ,
         \data_i[7][26] , \data_i[7][25] , \data_i[7][24] , \data_i[7][23] ,
         \data_i[7][22] , \data_i[7][21] , \data_i[7][20] , \data_i[7][19] ,
         \data_i[7][18] , \data_i[7][17] , \data_i[7][16] , \data_i[7][15] ,
         \data_i[7][14] , \data_i[7][13] , \data_i[7][12] , \data_i[7][11] ,
         \data_i[7][10] , \data_i[7][9] , \data_i[7][8] , \data_i[7][7] ,
         \data_i[7][6] , \data_i[7][5] , \data_i[7][4] , \data_i[7][3] ,
         \data_i[7][2] , \data_i[7][1] , \data_i[7][0] , \data_i[6][31] ,
         \data_i[6][30] , \data_i[6][29] , \data_i[6][28] , \data_i[6][27] ,
         \data_i[6][26] , \data_i[6][25] , \data_i[6][24] , \data_i[6][23] ,
         \data_i[6][22] , \data_i[6][21] , \data_i[6][20] , \data_i[6][19] ,
         \data_i[6][18] , \data_i[6][17] , \data_i[6][16] , \data_i[6][15] ,
         \data_i[6][14] , \data_i[6][13] , \data_i[6][12] , \data_i[6][11] ,
         \data_i[6][10] , \data_i[6][9] , \data_i[6][8] , \data_i[6][7] ,
         \data_i[6][6] , \data_i[6][5] , \data_i[6][4] , \data_i[6][3] ,
         \data_i[6][2] , \data_i[6][1] , \data_i[6][0] , \data_i[5][31] ,
         \data_i[5][30] , \data_i[5][29] , \data_i[5][28] , \data_i[5][27] ,
         \data_i[5][26] , \data_i[5][25] , \data_i[5][24] , \data_i[5][23] ,
         \data_i[5][22] , \data_i[5][21] , \data_i[5][20] , \data_i[5][19] ,
         \data_i[5][18] , \data_i[5][17] , \data_i[5][16] , \data_i[5][15] ,
         \data_i[5][14] , \data_i[5][13] , \data_i[5][12] , \data_i[5][11] ,
         \data_i[5][10] , \data_i[5][9] , \data_i[5][8] , \data_i[5][7] ,
         \data_i[5][6] , \data_i[5][5] , \data_i[5][4] , \data_i[5][3] ,
         \data_i[5][2] , \data_i[5][1] , \data_i[5][0] , \data_i[4][31] ,
         \data_i[4][30] , \data_i[4][29] , \data_i[4][28] , \data_i[4][27] ,
         \data_i[4][26] , \data_i[4][25] , \data_i[4][24] , \data_i[4][23] ,
         \data_i[4][22] , \data_i[4][21] , \data_i[4][20] , \data_i[4][19] ,
         \data_i[4][18] , \data_i[4][17] , \data_i[4][16] , \data_i[4][15] ,
         \data_i[4][14] , \data_i[4][13] , \data_i[4][12] , \data_i[4][11] ,
         \data_i[4][10] , \data_i[4][9] , \data_i[4][8] , \data_i[4][7] ,
         \data_i[4][6] , \data_i[4][5] , \data_i[4][4] , \data_i[4][3] ,
         \data_i[4][2] , \data_i[4][1] , \data_i[4][0] , \data_i[3][31] ,
         \data_i[3][30] , \data_i[3][29] , \data_i[3][28] , \data_i[3][27] ,
         \data_i[3][26] , \data_i[3][25] , \data_i[3][24] , \data_i[3][23] ,
         \data_i[3][22] , \data_i[3][21] , \data_i[3][20] , \data_i[3][19] ,
         \data_i[3][18] , \data_i[3][17] , \data_i[3][16] , \data_i[3][15] ,
         \data_i[3][14] , \data_i[3][13] , \data_i[3][12] , \data_i[3][11] ,
         \data_i[3][10] , \data_i[3][9] , \data_i[3][8] , \data_i[3][7] ,
         \data_i[3][6] , \data_i[3][5] , \data_i[3][4] , \data_i[3][3] ,
         \data_i[3][2] , \data_i[3][1] , \data_i[3][0] , \data_i[2][31] ,
         \data_i[2][30] , \data_i[2][29] , \data_i[2][28] , \data_i[2][27] ,
         \data_i[2][26] , \data_i[2][25] , \data_i[2][24] , \data_i[2][23] ,
         \data_i[2][22] , \data_i[2][21] , \data_i[2][20] , \data_i[2][19] ,
         \data_i[2][18] , \data_i[2][17] , \data_i[2][16] , \data_i[2][15] ,
         \data_i[2][14] , \data_i[2][13] , \data_i[2][12] , \data_i[2][11] ,
         \data_i[2][10] , \data_i[2][9] , \data_i[2][8] , \data_i[2][7] ,
         \data_i[2][6] , \data_i[2][5] , \data_i[2][4] , \data_i[2][3] ,
         \data_i[2][2] , \data_i[2][1] , \data_i[2][0] , \data_i[1][31] ,
         \data_i[1][30] , \data_i[1][29] , \data_i[1][28] , \data_i[1][27] ,
         \data_i[1][26] , \data_i[1][25] , \data_i[1][24] , \data_i[1][23] ,
         \data_i[1][22] , \data_i[1][21] , \data_i[1][20] , \data_i[1][19] ,
         \data_i[1][18] , \data_i[1][17] , \data_i[1][16] , \data_i[1][15] ,
         \data_i[1][14] , \data_i[1][13] , \data_i[1][12] , \data_i[1][11] ,
         \data_i[1][10] , \data_i[1][9] , \data_i[1][8] , \data_i[1][7] ,
         \data_i[1][6] , \data_i[1][5] , \data_i[1][4] , \data_i[1][3] ,
         \data_i[1][2] , \data_i[1][1] , \data_i[1][0] , \data_i[0][31] ,
         \data_i[0][30] , \data_i[0][29] , \data_i[0][28] , \data_i[0][27] ,
         \data_i[0][26] , \data_i[0][25] , \data_i[0][24] , \data_i[0][23] ,
         \data_i[0][22] , \data_i[0][21] , \data_i[0][20] , \data_i[0][19] ,
         \data_i[0][18] , \data_i[0][17] , \data_i[0][16] , \data_i[0][15] ,
         \data_i[0][14] , \data_i[0][13] , \data_i[0][12] , \data_i[0][11] ,
         \data_i[0][10] , \data_i[0][9] , \data_i[0][8] , \data_i[0][7] ,
         \data_i[0][6] , \data_i[0][5] , \data_i[0][4] , \data_i[0][3] ,
         \data_i[0][2] , \data_i[0][1] , \data_i[0][0] ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688;

  AND2X1_RVT U1 ( .A1(n24), .A2(n27), .Y(n675) );
  AND2X1_RVT U2 ( .A1(n24), .A2(n26), .Y(n676) );
  AND2X1_RVT U3 ( .A1(n23), .A2(n26), .Y(n673) );
  AND2X1_RVT U4 ( .A1(n18), .A2(n27), .Y(n667) );
  AND2X1_RVT U5 ( .A1(n18), .A2(n26), .Y(n668) );
  AND2X1_RVT U6 ( .A1(n17), .A2(n27), .Y(n663) );
  AND2X1_RVT U7 ( .A1(n17), .A2(n26), .Y(n664) );
  AND2X1_RVT U8 ( .A1(n16), .A2(n26), .Y(n661) );
  AND2X1_RVT U9 ( .A1(n16), .A2(n27), .Y(n662) );
  AND2X1_RVT U10 ( .A1(select_i[4]), .A2(n15), .Y(n27) );
  AND2X1_RVT U11 ( .A1(n10), .A2(n24), .Y(n651) );
  AND2X1_RVT U12 ( .A1(n9), .A2(n24), .Y(n652) );
  AND2X1_RVT U13 ( .A1(n9), .A2(n23), .Y(n649) );
  AND2X1_RVT U14 ( .A1(n10), .A2(n23), .Y(n650) );
  AND2X1_RVT U15 ( .A1(n10), .A2(n18), .Y(n643) );
  AND2X1_RVT U16 ( .A1(n9), .A2(n18), .Y(n644) );
  AND2X1_RVT U17 ( .A1(n10), .A2(n17), .Y(n639) );
  AND2X1_RVT U18 ( .A1(n9), .A2(n17), .Y(n640) );
  AND2X1_RVT U19 ( .A1(n16), .A2(n9), .Y(n637) );
  AND2X1_RVT U20 ( .A1(select_i[0]), .A2(n1), .Y(n9) );
  AND2X1_RVT U21 ( .A1(n10), .A2(n16), .Y(n638) );
  AND2X1_RVT U22 ( .A1(n1), .A2(n15), .Y(n10) );
  AND2X1_RVT U23 ( .A1(n28), .A2(n27), .Y(n679) );
  AND2X1_RVT U24 ( .A1(n28), .A2(n26), .Y(n680) );
  AND2X1_RVT U25 ( .A1(n25), .A2(n26), .Y(n677) );
  AND2X1_RVT U26 ( .A1(n25), .A2(n27), .Y(n678) );
  AND2X1_RVT U27 ( .A1(n23), .A2(n27), .Y(n674) );
  AND2X1_RVT U28 ( .A1(n10), .A2(n28), .Y(n655) );
  AND2X1_RVT U29 ( .A1(n9), .A2(n28), .Y(n656) );
  AND2X1_RVT U30 ( .A1(n9), .A2(n25), .Y(n653) );
  AND2X1_RVT U31 ( .A1(n10), .A2(n25), .Y(n654) );
  INVX1_RVT U32 ( .A(select_i[2]), .Y(n6) );
  AND2X1_RVT U33 ( .A1(select_i[4]), .A2(select_i[0]), .Y(n26) );
  INVX1_RVT U34 ( .A(select_i[1]), .Y(n8) );
  INVX1_RVT U35 ( .A(select_i[3]), .Y(n7) );
  INVX1_RVT U36 ( .A(select_i[0]), .Y(n15) );
  AND3X1_RVT U37 ( .A1(n6), .A2(n8), .A3(n7), .Y(n24) );
  AND3X1_RVT U38 ( .A1(select_i[1]), .A2(n6), .A3(n7), .Y(n23) );
  AND3X1_RVT U39 ( .A1(select_i[2]), .A2(select_i[3]), .A3(n8), .Y(n18) );
  AND3X1_RVT U40 ( .A1(select_i[3]), .A2(n6), .A3(n8), .Y(n17) );
  AND3X1_RVT U41 ( .A1(select_i[1]), .A2(select_i[3]), .A3(n6), .Y(n16) );
  INVX1_RVT U42 ( .A(select_i[4]), .Y(n1) );
  AND3X1_RVT U43 ( .A1(select_i[2]), .A2(n8), .A3(n7), .Y(n28) );
  AND3X1_RVT U44 ( .A1(select_i[1]), .A2(select_i[2]), .A3(n7), .Y(n25) );
  NAND4X0_RVT U45 ( .A1(n356), .A2(n355), .A3(n354), .A4(n353), .Y(data_o[24])
         );
  NAND4X0_RVT U46 ( .A1(n396), .A2(n395), .A3(n394), .A4(n393), .Y(data_o[26])
         );
  NAND4X0_RVT U47 ( .A1(n376), .A2(n375), .A3(n374), .A4(n373), .Y(data_o[25])
         );
  NAND4X0_RVT U48 ( .A1(n436), .A2(n435), .A3(n434), .A4(n433), .Y(data_o[28])
         );
  NAND4X0_RVT U49 ( .A1(n456), .A2(n455), .A3(n454), .A4(n453), .Y(data_o[29])
         );
  NAND4X0_RVT U50 ( .A1(n36), .A2(n35), .A3(n34), .A4(n33), .Y(data_o[0]) );
  NAND4X0_RVT U51 ( .A1(n256), .A2(n255), .A3(n254), .A4(n253), .Y(data_o[1])
         );
  NAND4X0_RVT U52 ( .A1(n416), .A2(n415), .A3(n414), .A4(n413), .Y(data_o[27])
         );
  NAND4X0_RVT U53 ( .A1(n536), .A2(n535), .A3(n534), .A4(n533), .Y(data_o[3])
         );
  NAND4X0_RVT U54 ( .A1(n556), .A2(n555), .A3(n554), .A4(n553), .Y(data_o[4])
         );
  NAND4X0_RVT U55 ( .A1(n576), .A2(n575), .A3(n574), .A4(n573), .Y(data_o[5])
         );
  NAND4X0_RVT U56 ( .A1(n596), .A2(n595), .A3(n594), .A4(n593), .Y(data_o[6])
         );
  NAND4X0_RVT U57 ( .A1(n616), .A2(n615), .A3(n614), .A4(n613), .Y(data_o[7])
         );
  NAND4X0_RVT U58 ( .A1(n636), .A2(n635), .A3(n634), .A4(n633), .Y(data_o[8])
         );
  NAND4X0_RVT U59 ( .A1(n688), .A2(n687), .A3(n686), .A4(n685), .Y(data_o[9])
         );
  NAND4X0_RVT U60 ( .A1(n56), .A2(n55), .A3(n54), .A4(n53), .Y(data_o[10]) );
  NAND4X0_RVT U61 ( .A1(n76), .A2(n75), .A3(n74), .A4(n73), .Y(data_o[11]) );
  NAND4X0_RVT U62 ( .A1(n96), .A2(n95), .A3(n94), .A4(n93), .Y(data_o[12]) );
  NAND4X0_RVT U63 ( .A1(n116), .A2(n115), .A3(n114), .A4(n113), .Y(data_o[13])
         );
  NAND4X0_RVT U64 ( .A1(n136), .A2(n135), .A3(n134), .A4(n133), .Y(data_o[14])
         );
  NAND4X0_RVT U65 ( .A1(n156), .A2(n155), .A3(n154), .A4(n153), .Y(data_o[15])
         );
  NAND4X0_RVT U66 ( .A1(n176), .A2(n175), .A3(n174), .A4(n173), .Y(data_o[16])
         );
  NAND4X0_RVT U67 ( .A1(n196), .A2(n195), .A3(n194), .A4(n193), .Y(data_o[17])
         );
  NAND4X0_RVT U68 ( .A1(n216), .A2(n215), .A3(n214), .A4(n213), .Y(data_o[18])
         );
  NAND4X0_RVT U69 ( .A1(n236), .A2(n235), .A3(n234), .A4(n233), .Y(data_o[19])
         );
  NAND4X0_RVT U70 ( .A1(n276), .A2(n275), .A3(n274), .A4(n273), .Y(data_o[20])
         );
  NAND4X0_RVT U71 ( .A1(n296), .A2(n295), .A3(n294), .A4(n293), .Y(data_o[21])
         );
  NAND4X0_RVT U72 ( .A1(n316), .A2(n315), .A3(n314), .A4(n313), .Y(data_o[22])
         );
  NAND4X0_RVT U73 ( .A1(n336), .A2(n335), .A3(n334), .A4(n333), .Y(data_o[23])
         );
  NAND4X0_RVT U74 ( .A1(n516), .A2(n515), .A3(n514), .A4(n513), .Y(data_o[31])
         );
  NAND4X0_RVT U75 ( .A1(n496), .A2(n495), .A3(n494), .A4(n493), .Y(data_o[30])
         );
  NAND4X0_RVT U76 ( .A1(n476), .A2(n475), .A3(n474), .A4(n473), .Y(data_o[2])
         );
  NOR4X1_RVT U77 ( .A1(n352), .A2(n351), .A3(n350), .A4(n349), .Y(n353) );
  NOR4X1_RVT U78 ( .A1(n348), .A2(n347), .A3(n346), .A4(n345), .Y(n354) );
  NOR4X1_RVT U79 ( .A1(n344), .A2(n343), .A3(n342), .A4(n341), .Y(n355) );
  NOR4X1_RVT U80 ( .A1(n340), .A2(n339), .A3(n338), .A4(n337), .Y(n356) );
  NOR4X1_RVT U81 ( .A1(n392), .A2(n391), .A3(n390), .A4(n389), .Y(n393) );
  NOR4X1_RVT U82 ( .A1(n388), .A2(n387), .A3(n386), .A4(n385), .Y(n394) );
  NOR4X1_RVT U83 ( .A1(n384), .A2(n383), .A3(n382), .A4(n381), .Y(n395) );
  NOR4X1_RVT U84 ( .A1(n380), .A2(n379), .A3(n378), .A4(n377), .Y(n396) );
  NOR4X1_RVT U85 ( .A1(n372), .A2(n371), .A3(n370), .A4(n369), .Y(n373) );
  NOR4X1_RVT U86 ( .A1(n368), .A2(n367), .A3(n366), .A4(n365), .Y(n374) );
  NOR4X1_RVT U87 ( .A1(n364), .A2(n363), .A3(n362), .A4(n361), .Y(n375) );
  NOR4X1_RVT U88 ( .A1(n360), .A2(n359), .A3(n358), .A4(n357), .Y(n376) );
  NOR4X1_RVT U89 ( .A1(n432), .A2(n431), .A3(n430), .A4(n429), .Y(n433) );
  NOR4X1_RVT U90 ( .A1(n428), .A2(n427), .A3(n426), .A4(n425), .Y(n434) );
  NOR4X1_RVT U91 ( .A1(n424), .A2(n423), .A3(n422), .A4(n421), .Y(n435) );
  NOR4X1_RVT U92 ( .A1(n420), .A2(n419), .A3(n418), .A4(n417), .Y(n436) );
  NOR4X1_RVT U93 ( .A1(n452), .A2(n451), .A3(n450), .A4(n449), .Y(n453) );
  NOR4X1_RVT U94 ( .A1(n448), .A2(n447), .A3(n446), .A4(n445), .Y(n454) );
  NOR4X1_RVT U95 ( .A1(n444), .A2(n443), .A3(n442), .A4(n441), .Y(n455) );
  NOR4X1_RVT U96 ( .A1(n440), .A2(n439), .A3(n438), .A4(n437), .Y(n456) );
  NOR4X1_RVT U97 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .Y(n33) );
  NOR4X1_RVT U98 ( .A1(n22), .A2(n21), .A3(n20), .A4(n19), .Y(n34) );
  NOR4X1_RVT U99 ( .A1(n14), .A2(n13), .A3(n12), .A4(n11), .Y(n35) );
  NOR4X1_RVT U100 ( .A1(n5), .A2(n4), .A3(n3), .A4(n2), .Y(n36) );
  NOR4X1_RVT U101 ( .A1(n252), .A2(n251), .A3(n250), .A4(n249), .Y(n253) );
  NOR4X1_RVT U102 ( .A1(n248), .A2(n247), .A3(n246), .A4(n245), .Y(n254) );
  NOR4X1_RVT U103 ( .A1(n244), .A2(n243), .A3(n242), .A4(n241), .Y(n255) );
  NOR4X1_RVT U104 ( .A1(n240), .A2(n239), .A3(n238), .A4(n237), .Y(n256) );
  NOR4X1_RVT U105 ( .A1(n412), .A2(n411), .A3(n410), .A4(n409), .Y(n413) );
  NOR4X1_RVT U106 ( .A1(n408), .A2(n407), .A3(n406), .A4(n405), .Y(n414) );
  NOR4X1_RVT U107 ( .A1(n404), .A2(n403), .A3(n402), .A4(n401), .Y(n415) );
  NOR4X1_RVT U108 ( .A1(n400), .A2(n399), .A3(n398), .A4(n397), .Y(n416) );
  NOR4X1_RVT U109 ( .A1(n532), .A2(n531), .A3(n530), .A4(n529), .Y(n533) );
  NOR4X1_RVT U110 ( .A1(n528), .A2(n527), .A3(n526), .A4(n525), .Y(n534) );
  NOR4X1_RVT U111 ( .A1(n524), .A2(n523), .A3(n522), .A4(n521), .Y(n535) );
  NOR4X1_RVT U112 ( .A1(n520), .A2(n519), .A3(n518), .A4(n517), .Y(n536) );
  NOR4X1_RVT U113 ( .A1(n552), .A2(n551), .A3(n550), .A4(n549), .Y(n553) );
  NOR4X1_RVT U114 ( .A1(n548), .A2(n547), .A3(n546), .A4(n545), .Y(n554) );
  NOR4X1_RVT U115 ( .A1(n544), .A2(n543), .A3(n542), .A4(n541), .Y(n555) );
  NOR4X1_RVT U116 ( .A1(n540), .A2(n539), .A3(n538), .A4(n537), .Y(n556) );
  NOR4X1_RVT U117 ( .A1(n572), .A2(n571), .A3(n570), .A4(n569), .Y(n573) );
  NOR4X1_RVT U118 ( .A1(n568), .A2(n567), .A3(n566), .A4(n565), .Y(n574) );
  NOR4X1_RVT U119 ( .A1(n564), .A2(n563), .A3(n562), .A4(n561), .Y(n575) );
  NOR4X1_RVT U120 ( .A1(n560), .A2(n559), .A3(n558), .A4(n557), .Y(n576) );
  NOR4X1_RVT U121 ( .A1(n592), .A2(n591), .A3(n590), .A4(n589), .Y(n593) );
  NOR4X1_RVT U122 ( .A1(n588), .A2(n587), .A3(n586), .A4(n585), .Y(n594) );
  NOR4X1_RVT U123 ( .A1(n584), .A2(n583), .A3(n582), .A4(n581), .Y(n595) );
  NOR4X1_RVT U124 ( .A1(n580), .A2(n579), .A3(n578), .A4(n577), .Y(n596) );
  NOR4X1_RVT U125 ( .A1(n612), .A2(n611), .A3(n610), .A4(n609), .Y(n613) );
  NOR4X1_RVT U126 ( .A1(n608), .A2(n607), .A3(n606), .A4(n605), .Y(n614) );
  NOR4X1_RVT U127 ( .A1(n604), .A2(n603), .A3(n602), .A4(n601), .Y(n615) );
  NOR4X1_RVT U128 ( .A1(n600), .A2(n599), .A3(n598), .A4(n597), .Y(n616) );
  NOR4X1_RVT U129 ( .A1(n632), .A2(n631), .A3(n630), .A4(n629), .Y(n633) );
  NOR4X1_RVT U130 ( .A1(n628), .A2(n627), .A3(n626), .A4(n625), .Y(n634) );
  NOR4X1_RVT U131 ( .A1(n624), .A2(n623), .A3(n622), .A4(n621), .Y(n635) );
  NOR4X1_RVT U132 ( .A1(n620), .A2(n619), .A3(n618), .A4(n617), .Y(n636) );
  NOR4X1_RVT U133 ( .A1(n684), .A2(n683), .A3(n682), .A4(n681), .Y(n685) );
  NOR4X1_RVT U134 ( .A1(n672), .A2(n671), .A3(n670), .A4(n669), .Y(n686) );
  NOR4X1_RVT U135 ( .A1(n660), .A2(n659), .A3(n658), .A4(n657), .Y(n687) );
  NOR4X1_RVT U136 ( .A1(n648), .A2(n647), .A3(n646), .A4(n645), .Y(n688) );
  NOR4X1_RVT U137 ( .A1(n52), .A2(n51), .A3(n50), .A4(n49), .Y(n53) );
  NOR4X1_RVT U138 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .Y(n54) );
  NOR4X1_RVT U139 ( .A1(n44), .A2(n43), .A3(n42), .A4(n41), .Y(n55) );
  NOR4X1_RVT U140 ( .A1(n40), .A2(n39), .A3(n38), .A4(n37), .Y(n56) );
  NOR4X1_RVT U141 ( .A1(n72), .A2(n71), .A3(n70), .A4(n69), .Y(n73) );
  NOR4X1_RVT U142 ( .A1(n68), .A2(n67), .A3(n66), .A4(n65), .Y(n74) );
  NOR4X1_RVT U143 ( .A1(n64), .A2(n63), .A3(n62), .A4(n61), .Y(n75) );
  NOR4X1_RVT U144 ( .A1(n60), .A2(n59), .A3(n58), .A4(n57), .Y(n76) );
  NOR4X1_RVT U145 ( .A1(n92), .A2(n91), .A3(n90), .A4(n89), .Y(n93) );
  NOR4X1_RVT U146 ( .A1(n88), .A2(n87), .A3(n86), .A4(n85), .Y(n94) );
  NOR4X1_RVT U147 ( .A1(n84), .A2(n83), .A3(n82), .A4(n81), .Y(n95) );
  NOR4X1_RVT U148 ( .A1(n80), .A2(n79), .A3(n78), .A4(n77), .Y(n96) );
  NOR4X1_RVT U149 ( .A1(n112), .A2(n111), .A3(n110), .A4(n109), .Y(n113) );
  NOR4X1_RVT U150 ( .A1(n108), .A2(n107), .A3(n106), .A4(n105), .Y(n114) );
  NOR4X1_RVT U151 ( .A1(n104), .A2(n103), .A3(n102), .A4(n101), .Y(n115) );
  NOR4X1_RVT U152 ( .A1(n100), .A2(n99), .A3(n98), .A4(n97), .Y(n116) );
  NOR4X1_RVT U153 ( .A1(n132), .A2(n131), .A3(n130), .A4(n129), .Y(n133) );
  NOR4X1_RVT U154 ( .A1(n128), .A2(n127), .A3(n126), .A4(n125), .Y(n134) );
  NOR4X1_RVT U155 ( .A1(n124), .A2(n123), .A3(n122), .A4(n121), .Y(n135) );
  NOR4X1_RVT U156 ( .A1(n120), .A2(n119), .A3(n118), .A4(n117), .Y(n136) );
  NOR4X1_RVT U157 ( .A1(n152), .A2(n151), .A3(n150), .A4(n149), .Y(n153) );
  NOR4X1_RVT U158 ( .A1(n148), .A2(n147), .A3(n146), .A4(n145), .Y(n154) );
  NOR4X1_RVT U159 ( .A1(n144), .A2(n143), .A3(n142), .A4(n141), .Y(n155) );
  NOR4X1_RVT U160 ( .A1(n140), .A2(n139), .A3(n138), .A4(n137), .Y(n156) );
  NOR4X1_RVT U161 ( .A1(n172), .A2(n171), .A3(n170), .A4(n169), .Y(n173) );
  NOR4X1_RVT U162 ( .A1(n168), .A2(n167), .A3(n166), .A4(n165), .Y(n174) );
  NOR4X1_RVT U163 ( .A1(n164), .A2(n163), .A3(n162), .A4(n161), .Y(n175) );
  NOR4X1_RVT U164 ( .A1(n160), .A2(n159), .A3(n158), .A4(n157), .Y(n176) );
  NOR4X1_RVT U165 ( .A1(n192), .A2(n191), .A3(n190), .A4(n189), .Y(n193) );
  NOR4X1_RVT U166 ( .A1(n188), .A2(n187), .A3(n186), .A4(n185), .Y(n194) );
  NOR4X1_RVT U167 ( .A1(n184), .A2(n183), .A3(n182), .A4(n181), .Y(n195) );
  NOR4X1_RVT U168 ( .A1(n180), .A2(n179), .A3(n178), .A4(n177), .Y(n196) );
  NOR4X1_RVT U169 ( .A1(n212), .A2(n211), .A3(n210), .A4(n209), .Y(n213) );
  NOR4X1_RVT U170 ( .A1(n208), .A2(n207), .A3(n206), .A4(n205), .Y(n214) );
  NOR4X1_RVT U171 ( .A1(n204), .A2(n203), .A3(n202), .A4(n201), .Y(n215) );
  NOR4X1_RVT U172 ( .A1(n200), .A2(n199), .A3(n198), .A4(n197), .Y(n216) );
  NOR4X1_RVT U173 ( .A1(n232), .A2(n231), .A3(n230), .A4(n229), .Y(n233) );
  NOR4X1_RVT U174 ( .A1(n228), .A2(n227), .A3(n226), .A4(n225), .Y(n234) );
  NOR4X1_RVT U175 ( .A1(n224), .A2(n223), .A3(n222), .A4(n221), .Y(n235) );
  NOR4X1_RVT U176 ( .A1(n220), .A2(n219), .A3(n218), .A4(n217), .Y(n236) );
  NOR4X1_RVT U177 ( .A1(n272), .A2(n271), .A3(n270), .A4(n269), .Y(n273) );
  NOR4X1_RVT U178 ( .A1(n268), .A2(n267), .A3(n266), .A4(n265), .Y(n274) );
  NOR4X1_RVT U179 ( .A1(n264), .A2(n263), .A3(n262), .A4(n261), .Y(n275) );
  NOR4X1_RVT U180 ( .A1(n260), .A2(n259), .A3(n258), .A4(n257), .Y(n276) );
  NOR4X1_RVT U181 ( .A1(n292), .A2(n291), .A3(n290), .A4(n289), .Y(n293) );
  NOR4X1_RVT U182 ( .A1(n288), .A2(n287), .A3(n286), .A4(n285), .Y(n294) );
  NOR4X1_RVT U183 ( .A1(n284), .A2(n283), .A3(n282), .A4(n281), .Y(n295) );
  NOR4X1_RVT U184 ( .A1(n280), .A2(n279), .A3(n278), .A4(n277), .Y(n296) );
  NOR4X1_RVT U185 ( .A1(n312), .A2(n311), .A3(n310), .A4(n309), .Y(n313) );
  NOR4X1_RVT U186 ( .A1(n308), .A2(n307), .A3(n306), .A4(n305), .Y(n314) );
  NOR4X1_RVT U187 ( .A1(n304), .A2(n303), .A3(n302), .A4(n301), .Y(n315) );
  NOR4X1_RVT U188 ( .A1(n300), .A2(n299), .A3(n298), .A4(n297), .Y(n316) );
  NOR4X1_RVT U189 ( .A1(n332), .A2(n331), .A3(n330), .A4(n329), .Y(n333) );
  NOR4X1_RVT U190 ( .A1(n328), .A2(n327), .A3(n326), .A4(n325), .Y(n334) );
  NOR4X1_RVT U191 ( .A1(n324), .A2(n323), .A3(n322), .A4(n321), .Y(n335) );
  NOR4X1_RVT U192 ( .A1(n320), .A2(n319), .A3(n318), .A4(n317), .Y(n336) );
  NOR4X1_RVT U193 ( .A1(n512), .A2(n511), .A3(n510), .A4(n509), .Y(n513) );
  NOR4X1_RVT U194 ( .A1(n508), .A2(n507), .A3(n506), .A4(n505), .Y(n514) );
  NOR4X1_RVT U195 ( .A1(n504), .A2(n503), .A3(n502), .A4(n501), .Y(n515) );
  NOR4X1_RVT U196 ( .A1(n500), .A2(n499), .A3(n498), .A4(n497), .Y(n516) );
  NOR4X1_RVT U197 ( .A1(n492), .A2(n491), .A3(n490), .A4(n489), .Y(n493) );
  NOR4X1_RVT U198 ( .A1(n488), .A2(n487), .A3(n486), .A4(n485), .Y(n494) );
  NOR4X1_RVT U199 ( .A1(n484), .A2(n483), .A3(n482), .A4(n481), .Y(n495) );
  NOR4X1_RVT U200 ( .A1(n480), .A2(n479), .A3(n478), .A4(n477), .Y(n496) );
  NOR4X1_RVT U201 ( .A1(n472), .A2(n471), .A3(n470), .A4(n469), .Y(n473) );
  NOR4X1_RVT U202 ( .A1(n468), .A2(n467), .A3(n466), .A4(n465), .Y(n474) );
  AND4X1_RVT U203 ( .A1(select_i[2]), .A2(select_i[1]), .A3(select_i[3]), .A4(
        n26), .Y(n665) );
  AND4X1_RVT U204 ( .A1(select_i[2]), .A2(select_i[1]), .A3(select_i[3]), .A4(
        n27), .Y(n666) );
  NOR4X1_RVT U205 ( .A1(n464), .A2(n463), .A3(n462), .A4(n461), .Y(n475) );
  NOR4X1_RVT U206 ( .A1(n460), .A2(n459), .A3(n458), .A4(n457), .Y(n476) );
  AND4X1_RVT U207 ( .A1(select_i[2]), .A2(select_i[1]), .A3(select_i[3]), .A4(
        n9), .Y(n641) );
  AND4X1_RVT U208 ( .A1(n10), .A2(select_i[2]), .A3(select_i[1]), .A4(
        select_i[3]), .Y(n642) );
  AO22X1_RVT U209 ( .A1(n638), .A2(\data_i[10][0] ), .A3(n637), .A4(
        \data_i[11][0] ), .Y(n5) );
  AO22X1_RVT U210 ( .A1(n640), .A2(\data_i[9][0] ), .A3(n639), .A4(
        \data_i[8][0] ), .Y(n4) );
  AO22X1_RVT U211 ( .A1(n642), .A2(\data_i[14][0] ), .A3(n641), .A4(
        \data_i[15][0] ), .Y(n3) );
  AO22X1_RVT U212 ( .A1(n644), .A2(\data_i[13][0] ), .A3(n643), .A4(
        \data_i[12][0] ), .Y(n2) );
  AO22X1_RVT U213 ( .A1(n650), .A2(\data_i[2][0] ), .A3(n649), .A4(
        \data_i[3][0] ), .Y(n14) );
  AO22X1_RVT U214 ( .A1(n652), .A2(\data_i[1][0] ), .A3(n651), .A4(
        \data_i[0][0] ), .Y(n13) );
  AO22X1_RVT U215 ( .A1(n654), .A2(\data_i[6][0] ), .A3(n653), .A4(
        \data_i[7][0] ), .Y(n12) );
  AO22X1_RVT U216 ( .A1(n656), .A2(\data_i[5][0] ), .A3(n655), .A4(
        \data_i[4][0] ), .Y(n11) );
  AO22X1_RVT U217 ( .A1(n662), .A2(\data_i[26][0] ), .A3(n661), .A4(
        \data_i[27][0] ), .Y(n22) );
  AO22X1_RVT U218 ( .A1(n664), .A2(\data_i[25][0] ), .A3(n663), .A4(
        \data_i[24][0] ), .Y(n21) );
  AO22X1_RVT U219 ( .A1(n666), .A2(\data_i[30][0] ), .A3(n665), .A4(
        \data_i[31][0] ), .Y(n20) );
  AO22X1_RVT U220 ( .A1(n668), .A2(\data_i[29][0] ), .A3(n667), .A4(
        \data_i[28][0] ), .Y(n19) );
  AO22X1_RVT U221 ( .A1(n674), .A2(\data_i[18][0] ), .A3(n673), .A4(
        \data_i[19][0] ), .Y(n32) );
  AO22X1_RVT U222 ( .A1(n676), .A2(\data_i[17][0] ), .A3(n675), .A4(
        \data_i[16][0] ), .Y(n31) );
  AO22X1_RVT U223 ( .A1(n678), .A2(\data_i[22][0] ), .A3(n677), .A4(
        \data_i[23][0] ), .Y(n30) );
  AO22X1_RVT U224 ( .A1(n680), .A2(\data_i[21][0] ), .A3(n679), .A4(
        \data_i[20][0] ), .Y(n29) );
  AO22X1_RVT U225 ( .A1(n638), .A2(\data_i[10][10] ), .A3(n637), .A4(
        \data_i[11][10] ), .Y(n40) );
  AO22X1_RVT U226 ( .A1(n640), .A2(\data_i[9][10] ), .A3(n639), .A4(
        \data_i[8][10] ), .Y(n39) );
  AO22X1_RVT U227 ( .A1(n642), .A2(\data_i[14][10] ), .A3(n641), .A4(
        \data_i[15][10] ), .Y(n38) );
  AO22X1_RVT U228 ( .A1(n644), .A2(\data_i[13][10] ), .A3(n643), .A4(
        \data_i[12][10] ), .Y(n37) );
  AO22X1_RVT U229 ( .A1(n650), .A2(\data_i[2][10] ), .A3(n649), .A4(
        \data_i[3][10] ), .Y(n44) );
  AO22X1_RVT U230 ( .A1(n652), .A2(\data_i[1][10] ), .A3(n651), .A4(
        \data_i[0][10] ), .Y(n43) );
  AO22X1_RVT U231 ( .A1(n654), .A2(\data_i[6][10] ), .A3(n653), .A4(
        \data_i[7][10] ), .Y(n42) );
  AO22X1_RVT U232 ( .A1(n656), .A2(\data_i[5][10] ), .A3(n655), .A4(
        \data_i[4][10] ), .Y(n41) );
  AO22X1_RVT U233 ( .A1(n662), .A2(\data_i[26][10] ), .A3(n661), .A4(
        \data_i[27][10] ), .Y(n48) );
  AO22X1_RVT U234 ( .A1(n664), .A2(\data_i[25][10] ), .A3(n663), .A4(
        \data_i[24][10] ), .Y(n47) );
  AO22X1_RVT U235 ( .A1(n666), .A2(\data_i[30][10] ), .A3(n665), .A4(
        \data_i[31][10] ), .Y(n46) );
  AO22X1_RVT U236 ( .A1(n668), .A2(\data_i[29][10] ), .A3(n667), .A4(
        \data_i[28][10] ), .Y(n45) );
  AO22X1_RVT U237 ( .A1(n674), .A2(\data_i[18][10] ), .A3(n673), .A4(
        \data_i[19][10] ), .Y(n52) );
  AO22X1_RVT U238 ( .A1(n676), .A2(\data_i[17][10] ), .A3(n675), .A4(
        \data_i[16][10] ), .Y(n51) );
  AO22X1_RVT U239 ( .A1(n678), .A2(\data_i[22][10] ), .A3(n677), .A4(
        \data_i[23][10] ), .Y(n50) );
  AO22X1_RVT U240 ( .A1(n680), .A2(\data_i[21][10] ), .A3(n679), .A4(
        \data_i[20][10] ), .Y(n49) );
  AO22X1_RVT U241 ( .A1(n638), .A2(\data_i[10][11] ), .A3(n637), .A4(
        \data_i[11][11] ), .Y(n60) );
  AO22X1_RVT U242 ( .A1(n640), .A2(\data_i[9][11] ), .A3(n639), .A4(
        \data_i[8][11] ), .Y(n59) );
  AO22X1_RVT U243 ( .A1(n642), .A2(\data_i[14][11] ), .A3(n641), .A4(
        \data_i[15][11] ), .Y(n58) );
  AO22X1_RVT U244 ( .A1(n644), .A2(\data_i[13][11] ), .A3(n643), .A4(
        \data_i[12][11] ), .Y(n57) );
  AO22X1_RVT U245 ( .A1(n650), .A2(\data_i[2][11] ), .A3(n649), .A4(
        \data_i[3][11] ), .Y(n64) );
  AO22X1_RVT U246 ( .A1(n652), .A2(\data_i[1][11] ), .A3(n651), .A4(
        \data_i[0][11] ), .Y(n63) );
  AO22X1_RVT U247 ( .A1(n654), .A2(\data_i[6][11] ), .A3(n653), .A4(
        \data_i[7][11] ), .Y(n62) );
  AO22X1_RVT U248 ( .A1(n656), .A2(\data_i[5][11] ), .A3(n655), .A4(
        \data_i[4][11] ), .Y(n61) );
  AO22X1_RVT U249 ( .A1(n662), .A2(\data_i[26][11] ), .A3(n661), .A4(
        \data_i[27][11] ), .Y(n68) );
  AO22X1_RVT U250 ( .A1(n664), .A2(\data_i[25][11] ), .A3(n663), .A4(
        \data_i[24][11] ), .Y(n67) );
  AO22X1_RVT U251 ( .A1(n666), .A2(\data_i[30][11] ), .A3(n665), .A4(
        \data_i[31][11] ), .Y(n66) );
  AO22X1_RVT U252 ( .A1(n668), .A2(\data_i[29][11] ), .A3(n667), .A4(
        \data_i[28][11] ), .Y(n65) );
  AO22X1_RVT U253 ( .A1(n674), .A2(\data_i[18][11] ), .A3(n673), .A4(
        \data_i[19][11] ), .Y(n72) );
  AO22X1_RVT U254 ( .A1(n676), .A2(\data_i[17][11] ), .A3(n675), .A4(
        \data_i[16][11] ), .Y(n71) );
  AO22X1_RVT U255 ( .A1(n678), .A2(\data_i[22][11] ), .A3(n677), .A4(
        \data_i[23][11] ), .Y(n70) );
  AO22X1_RVT U256 ( .A1(n680), .A2(\data_i[21][11] ), .A3(n679), .A4(
        \data_i[20][11] ), .Y(n69) );
  AO22X1_RVT U257 ( .A1(n638), .A2(\data_i[10][12] ), .A3(n637), .A4(
        \data_i[11][12] ), .Y(n80) );
  AO22X1_RVT U258 ( .A1(n640), .A2(\data_i[9][12] ), .A3(n639), .A4(
        \data_i[8][12] ), .Y(n79) );
  AO22X1_RVT U259 ( .A1(n642), .A2(\data_i[14][12] ), .A3(n641), .A4(
        \data_i[15][12] ), .Y(n78) );
  AO22X1_RVT U260 ( .A1(n644), .A2(\data_i[13][12] ), .A3(n643), .A4(
        \data_i[12][12] ), .Y(n77) );
  AO22X1_RVT U261 ( .A1(n650), .A2(\data_i[2][12] ), .A3(n649), .A4(
        \data_i[3][12] ), .Y(n84) );
  AO22X1_RVT U262 ( .A1(n652), .A2(\data_i[1][12] ), .A3(n651), .A4(
        \data_i[0][12] ), .Y(n83) );
  AO22X1_RVT U263 ( .A1(n654), .A2(\data_i[6][12] ), .A3(n653), .A4(
        \data_i[7][12] ), .Y(n82) );
  AO22X1_RVT U264 ( .A1(n656), .A2(\data_i[5][12] ), .A3(n655), .A4(
        \data_i[4][12] ), .Y(n81) );
  AO22X1_RVT U265 ( .A1(n662), .A2(\data_i[26][12] ), .A3(n661), .A4(
        \data_i[27][12] ), .Y(n88) );
  AO22X1_RVT U266 ( .A1(n664), .A2(\data_i[25][12] ), .A3(n663), .A4(
        \data_i[24][12] ), .Y(n87) );
  AO22X1_RVT U267 ( .A1(n666), .A2(\data_i[30][12] ), .A3(n665), .A4(
        \data_i[31][12] ), .Y(n86) );
  AO22X1_RVT U268 ( .A1(n668), .A2(\data_i[29][12] ), .A3(n667), .A4(
        \data_i[28][12] ), .Y(n85) );
  AO22X1_RVT U269 ( .A1(n674), .A2(\data_i[18][12] ), .A3(n673), .A4(
        \data_i[19][12] ), .Y(n92) );
  AO22X1_RVT U270 ( .A1(n676), .A2(\data_i[17][12] ), .A3(n675), .A4(
        \data_i[16][12] ), .Y(n91) );
  AO22X1_RVT U271 ( .A1(n678), .A2(\data_i[22][12] ), .A3(n677), .A4(
        \data_i[23][12] ), .Y(n90) );
  AO22X1_RVT U272 ( .A1(n680), .A2(\data_i[21][12] ), .A3(n679), .A4(
        \data_i[20][12] ), .Y(n89) );
  AO22X1_RVT U273 ( .A1(n638), .A2(\data_i[10][13] ), .A3(n637), .A4(
        \data_i[11][13] ), .Y(n100) );
  AO22X1_RVT U274 ( .A1(n640), .A2(\data_i[9][13] ), .A3(n639), .A4(
        \data_i[8][13] ), .Y(n99) );
  AO22X1_RVT U275 ( .A1(n642), .A2(\data_i[14][13] ), .A3(n641), .A4(
        \data_i[15][13] ), .Y(n98) );
  AO22X1_RVT U276 ( .A1(n644), .A2(\data_i[13][13] ), .A3(n643), .A4(
        \data_i[12][13] ), .Y(n97) );
  AO22X1_RVT U277 ( .A1(n650), .A2(\data_i[2][13] ), .A3(n649), .A4(
        \data_i[3][13] ), .Y(n104) );
  AO22X1_RVT U278 ( .A1(n652), .A2(\data_i[1][13] ), .A3(n651), .A4(
        \data_i[0][13] ), .Y(n103) );
  AO22X1_RVT U279 ( .A1(n654), .A2(\data_i[6][13] ), .A3(n653), .A4(
        \data_i[7][13] ), .Y(n102) );
  AO22X1_RVT U280 ( .A1(n656), .A2(\data_i[5][13] ), .A3(n655), .A4(
        \data_i[4][13] ), .Y(n101) );
  AO22X1_RVT U281 ( .A1(n662), .A2(\data_i[26][13] ), .A3(n661), .A4(
        \data_i[27][13] ), .Y(n108) );
  AO22X1_RVT U282 ( .A1(n664), .A2(\data_i[25][13] ), .A3(n663), .A4(
        \data_i[24][13] ), .Y(n107) );
  AO22X1_RVT U283 ( .A1(n666), .A2(\data_i[30][13] ), .A3(n665), .A4(
        \data_i[31][13] ), .Y(n106) );
  AO22X1_RVT U284 ( .A1(n668), .A2(\data_i[29][13] ), .A3(n667), .A4(
        \data_i[28][13] ), .Y(n105) );
  AO22X1_RVT U285 ( .A1(n674), .A2(\data_i[18][13] ), .A3(n673), .A4(
        \data_i[19][13] ), .Y(n112) );
  AO22X1_RVT U286 ( .A1(n676), .A2(\data_i[17][13] ), .A3(n675), .A4(
        \data_i[16][13] ), .Y(n111) );
  AO22X1_RVT U287 ( .A1(n678), .A2(\data_i[22][13] ), .A3(n677), .A4(
        \data_i[23][13] ), .Y(n110) );
  AO22X1_RVT U288 ( .A1(n680), .A2(\data_i[21][13] ), .A3(n679), .A4(
        \data_i[20][13] ), .Y(n109) );
  AO22X1_RVT U289 ( .A1(n638), .A2(\data_i[10][14] ), .A3(n637), .A4(
        \data_i[11][14] ), .Y(n120) );
  AO22X1_RVT U290 ( .A1(n640), .A2(\data_i[9][14] ), .A3(n639), .A4(
        \data_i[8][14] ), .Y(n119) );
  AO22X1_RVT U291 ( .A1(n642), .A2(\data_i[14][14] ), .A3(n641), .A4(
        \data_i[15][14] ), .Y(n118) );
  AO22X1_RVT U292 ( .A1(n644), .A2(\data_i[13][14] ), .A3(n643), .A4(
        \data_i[12][14] ), .Y(n117) );
  AO22X1_RVT U293 ( .A1(n650), .A2(\data_i[2][14] ), .A3(n649), .A4(
        \data_i[3][14] ), .Y(n124) );
  AO22X1_RVT U294 ( .A1(n652), .A2(\data_i[1][14] ), .A3(n651), .A4(
        \data_i[0][14] ), .Y(n123) );
  AO22X1_RVT U295 ( .A1(n654), .A2(\data_i[6][14] ), .A3(n653), .A4(
        \data_i[7][14] ), .Y(n122) );
  AO22X1_RVT U296 ( .A1(n656), .A2(\data_i[5][14] ), .A3(n655), .A4(
        \data_i[4][14] ), .Y(n121) );
  AO22X1_RVT U297 ( .A1(n662), .A2(\data_i[26][14] ), .A3(n661), .A4(
        \data_i[27][14] ), .Y(n128) );
  AO22X1_RVT U298 ( .A1(n664), .A2(\data_i[25][14] ), .A3(n663), .A4(
        \data_i[24][14] ), .Y(n127) );
  AO22X1_RVT U299 ( .A1(n666), .A2(\data_i[30][14] ), .A3(n665), .A4(
        \data_i[31][14] ), .Y(n126) );
  AO22X1_RVT U300 ( .A1(n668), .A2(\data_i[29][14] ), .A3(n667), .A4(
        \data_i[28][14] ), .Y(n125) );
  AO22X1_RVT U301 ( .A1(n674), .A2(\data_i[18][14] ), .A3(n673), .A4(
        \data_i[19][14] ), .Y(n132) );
  AO22X1_RVT U302 ( .A1(n676), .A2(\data_i[17][14] ), .A3(n675), .A4(
        \data_i[16][14] ), .Y(n131) );
  AO22X1_RVT U303 ( .A1(n678), .A2(\data_i[22][14] ), .A3(n677), .A4(
        \data_i[23][14] ), .Y(n130) );
  AO22X1_RVT U304 ( .A1(n680), .A2(\data_i[21][14] ), .A3(n679), .A4(
        \data_i[20][14] ), .Y(n129) );
  AO22X1_RVT U305 ( .A1(n638), .A2(\data_i[10][15] ), .A3(n637), .A4(
        \data_i[11][15] ), .Y(n140) );
  AO22X1_RVT U306 ( .A1(n640), .A2(\data_i[9][15] ), .A3(n639), .A4(
        \data_i[8][15] ), .Y(n139) );
  AO22X1_RVT U307 ( .A1(n642), .A2(\data_i[14][15] ), .A3(n641), .A4(
        \data_i[15][15] ), .Y(n138) );
  AO22X1_RVT U308 ( .A1(n644), .A2(\data_i[13][15] ), .A3(n643), .A4(
        \data_i[12][15] ), .Y(n137) );
  AO22X1_RVT U309 ( .A1(n650), .A2(\data_i[2][15] ), .A3(n649), .A4(
        \data_i[3][15] ), .Y(n144) );
  AO22X1_RVT U310 ( .A1(n652), .A2(\data_i[1][15] ), .A3(n651), .A4(
        \data_i[0][15] ), .Y(n143) );
  AO22X1_RVT U311 ( .A1(n654), .A2(\data_i[6][15] ), .A3(n653), .A4(
        \data_i[7][15] ), .Y(n142) );
  AO22X1_RVT U312 ( .A1(n656), .A2(\data_i[5][15] ), .A3(n655), .A4(
        \data_i[4][15] ), .Y(n141) );
  AO22X1_RVT U313 ( .A1(n662), .A2(\data_i[26][15] ), .A3(n661), .A4(
        \data_i[27][15] ), .Y(n148) );
  AO22X1_RVT U314 ( .A1(n664), .A2(\data_i[25][15] ), .A3(n663), .A4(
        \data_i[24][15] ), .Y(n147) );
  AO22X1_RVT U315 ( .A1(n666), .A2(\data_i[30][15] ), .A3(n665), .A4(
        \data_i[31][15] ), .Y(n146) );
  AO22X1_RVT U316 ( .A1(n668), .A2(\data_i[29][15] ), .A3(n667), .A4(
        \data_i[28][15] ), .Y(n145) );
  AO22X1_RVT U317 ( .A1(n674), .A2(\data_i[18][15] ), .A3(n673), .A4(
        \data_i[19][15] ), .Y(n152) );
  AO22X1_RVT U318 ( .A1(n676), .A2(\data_i[17][15] ), .A3(n675), .A4(
        \data_i[16][15] ), .Y(n151) );
  AO22X1_RVT U319 ( .A1(n678), .A2(\data_i[22][15] ), .A3(n677), .A4(
        \data_i[23][15] ), .Y(n150) );
  AO22X1_RVT U320 ( .A1(n680), .A2(\data_i[21][15] ), .A3(n679), .A4(
        \data_i[20][15] ), .Y(n149) );
  AO22X1_RVT U321 ( .A1(n638), .A2(\data_i[10][16] ), .A3(n637), .A4(
        \data_i[11][16] ), .Y(n160) );
  AO22X1_RVT U322 ( .A1(n640), .A2(\data_i[9][16] ), .A3(n639), .A4(
        \data_i[8][16] ), .Y(n159) );
  AO22X1_RVT U323 ( .A1(n642), .A2(\data_i[14][16] ), .A3(n641), .A4(
        \data_i[15][16] ), .Y(n158) );
  AO22X1_RVT U324 ( .A1(n644), .A2(\data_i[13][16] ), .A3(n643), .A4(
        \data_i[12][16] ), .Y(n157) );
  AO22X1_RVT U325 ( .A1(n650), .A2(\data_i[2][16] ), .A3(n649), .A4(
        \data_i[3][16] ), .Y(n164) );
  AO22X1_RVT U326 ( .A1(n652), .A2(\data_i[1][16] ), .A3(n651), .A4(
        \data_i[0][16] ), .Y(n163) );
  AO22X1_RVT U327 ( .A1(n654), .A2(\data_i[6][16] ), .A3(n653), .A4(
        \data_i[7][16] ), .Y(n162) );
  AO22X1_RVT U328 ( .A1(n656), .A2(\data_i[5][16] ), .A3(n655), .A4(
        \data_i[4][16] ), .Y(n161) );
  AO22X1_RVT U329 ( .A1(n662), .A2(\data_i[26][16] ), .A3(n661), .A4(
        \data_i[27][16] ), .Y(n168) );
  AO22X1_RVT U330 ( .A1(n664), .A2(\data_i[25][16] ), .A3(n663), .A4(
        \data_i[24][16] ), .Y(n167) );
  AO22X1_RVT U331 ( .A1(n666), .A2(\data_i[30][16] ), .A3(n665), .A4(
        \data_i[31][16] ), .Y(n166) );
  AO22X1_RVT U332 ( .A1(n668), .A2(\data_i[29][16] ), .A3(n667), .A4(
        \data_i[28][16] ), .Y(n165) );
  AO22X1_RVT U333 ( .A1(n674), .A2(\data_i[18][16] ), .A3(n673), .A4(
        \data_i[19][16] ), .Y(n172) );
  AO22X1_RVT U334 ( .A1(n676), .A2(\data_i[17][16] ), .A3(n675), .A4(
        \data_i[16][16] ), .Y(n171) );
  AO22X1_RVT U335 ( .A1(n678), .A2(\data_i[22][16] ), .A3(n677), .A4(
        \data_i[23][16] ), .Y(n170) );
  AO22X1_RVT U336 ( .A1(n680), .A2(\data_i[21][16] ), .A3(n679), .A4(
        \data_i[20][16] ), .Y(n169) );
  AO22X1_RVT U337 ( .A1(n638), .A2(\data_i[10][17] ), .A3(n637), .A4(
        \data_i[11][17] ), .Y(n180) );
  AO22X1_RVT U338 ( .A1(n640), .A2(\data_i[9][17] ), .A3(n639), .A4(
        \data_i[8][17] ), .Y(n179) );
  AO22X1_RVT U339 ( .A1(n642), .A2(\data_i[14][17] ), .A3(n641), .A4(
        \data_i[15][17] ), .Y(n178) );
  AO22X1_RVT U340 ( .A1(n644), .A2(\data_i[13][17] ), .A3(n643), .A4(
        \data_i[12][17] ), .Y(n177) );
  AO22X1_RVT U341 ( .A1(n650), .A2(\data_i[2][17] ), .A3(n649), .A4(
        \data_i[3][17] ), .Y(n184) );
  AO22X1_RVT U342 ( .A1(n652), .A2(\data_i[1][17] ), .A3(n651), .A4(
        \data_i[0][17] ), .Y(n183) );
  AO22X1_RVT U343 ( .A1(n654), .A2(\data_i[6][17] ), .A3(n653), .A4(
        \data_i[7][17] ), .Y(n182) );
  AO22X1_RVT U344 ( .A1(n656), .A2(\data_i[5][17] ), .A3(n655), .A4(
        \data_i[4][17] ), .Y(n181) );
  AO22X1_RVT U345 ( .A1(n662), .A2(\data_i[26][17] ), .A3(n661), .A4(
        \data_i[27][17] ), .Y(n188) );
  AO22X1_RVT U346 ( .A1(n664), .A2(\data_i[25][17] ), .A3(n663), .A4(
        \data_i[24][17] ), .Y(n187) );
  AO22X1_RVT U347 ( .A1(n666), .A2(\data_i[30][17] ), .A3(n665), .A4(
        \data_i[31][17] ), .Y(n186) );
  AO22X1_RVT U348 ( .A1(n668), .A2(\data_i[29][17] ), .A3(n667), .A4(
        \data_i[28][17] ), .Y(n185) );
  AO22X1_RVT U349 ( .A1(n674), .A2(\data_i[18][17] ), .A3(n673), .A4(
        \data_i[19][17] ), .Y(n192) );
  AO22X1_RVT U350 ( .A1(n676), .A2(\data_i[17][17] ), .A3(n675), .A4(
        \data_i[16][17] ), .Y(n191) );
  AO22X1_RVT U351 ( .A1(n678), .A2(\data_i[22][17] ), .A3(n677), .A4(
        \data_i[23][17] ), .Y(n190) );
  AO22X1_RVT U352 ( .A1(n680), .A2(\data_i[21][17] ), .A3(n679), .A4(
        \data_i[20][17] ), .Y(n189) );
  AO22X1_RVT U353 ( .A1(n638), .A2(\data_i[10][18] ), .A3(n637), .A4(
        \data_i[11][18] ), .Y(n200) );
  AO22X1_RVT U354 ( .A1(n640), .A2(\data_i[9][18] ), .A3(n639), .A4(
        \data_i[8][18] ), .Y(n199) );
  AO22X1_RVT U355 ( .A1(n642), .A2(\data_i[14][18] ), .A3(n641), .A4(
        \data_i[15][18] ), .Y(n198) );
  AO22X1_RVT U356 ( .A1(n644), .A2(\data_i[13][18] ), .A3(n643), .A4(
        \data_i[12][18] ), .Y(n197) );
  AO22X1_RVT U357 ( .A1(n650), .A2(\data_i[2][18] ), .A3(n649), .A4(
        \data_i[3][18] ), .Y(n204) );
  AO22X1_RVT U358 ( .A1(n652), .A2(\data_i[1][18] ), .A3(n651), .A4(
        \data_i[0][18] ), .Y(n203) );
  AO22X1_RVT U359 ( .A1(n654), .A2(\data_i[6][18] ), .A3(n653), .A4(
        \data_i[7][18] ), .Y(n202) );
  AO22X1_RVT U360 ( .A1(n656), .A2(\data_i[5][18] ), .A3(n655), .A4(
        \data_i[4][18] ), .Y(n201) );
  AO22X1_RVT U361 ( .A1(n662), .A2(\data_i[26][18] ), .A3(n661), .A4(
        \data_i[27][18] ), .Y(n208) );
  AO22X1_RVT U362 ( .A1(n664), .A2(\data_i[25][18] ), .A3(n663), .A4(
        \data_i[24][18] ), .Y(n207) );
  AO22X1_RVT U363 ( .A1(n666), .A2(\data_i[30][18] ), .A3(n665), .A4(
        \data_i[31][18] ), .Y(n206) );
  AO22X1_RVT U364 ( .A1(n668), .A2(\data_i[29][18] ), .A3(n667), .A4(
        \data_i[28][18] ), .Y(n205) );
  AO22X1_RVT U365 ( .A1(n674), .A2(\data_i[18][18] ), .A3(n673), .A4(
        \data_i[19][18] ), .Y(n212) );
  AO22X1_RVT U366 ( .A1(n676), .A2(\data_i[17][18] ), .A3(n675), .A4(
        \data_i[16][18] ), .Y(n211) );
  AO22X1_RVT U367 ( .A1(n678), .A2(\data_i[22][18] ), .A3(n677), .A4(
        \data_i[23][18] ), .Y(n210) );
  AO22X1_RVT U368 ( .A1(n680), .A2(\data_i[21][18] ), .A3(n679), .A4(
        \data_i[20][18] ), .Y(n209) );
  AO22X1_RVT U369 ( .A1(n638), .A2(\data_i[10][19] ), .A3(n637), .A4(
        \data_i[11][19] ), .Y(n220) );
  AO22X1_RVT U370 ( .A1(n640), .A2(\data_i[9][19] ), .A3(n639), .A4(
        \data_i[8][19] ), .Y(n219) );
  AO22X1_RVT U371 ( .A1(n642), .A2(\data_i[14][19] ), .A3(n641), .A4(
        \data_i[15][19] ), .Y(n218) );
  AO22X1_RVT U372 ( .A1(n644), .A2(\data_i[13][19] ), .A3(n643), .A4(
        \data_i[12][19] ), .Y(n217) );
  AO22X1_RVT U373 ( .A1(n650), .A2(\data_i[2][19] ), .A3(n649), .A4(
        \data_i[3][19] ), .Y(n224) );
  AO22X1_RVT U374 ( .A1(n652), .A2(\data_i[1][19] ), .A3(n651), .A4(
        \data_i[0][19] ), .Y(n223) );
  AO22X1_RVT U375 ( .A1(n654), .A2(\data_i[6][19] ), .A3(n653), .A4(
        \data_i[7][19] ), .Y(n222) );
  AO22X1_RVT U376 ( .A1(n656), .A2(\data_i[5][19] ), .A3(n655), .A4(
        \data_i[4][19] ), .Y(n221) );
  AO22X1_RVT U377 ( .A1(n662), .A2(\data_i[26][19] ), .A3(n661), .A4(
        \data_i[27][19] ), .Y(n228) );
  AO22X1_RVT U378 ( .A1(n664), .A2(\data_i[25][19] ), .A3(n663), .A4(
        \data_i[24][19] ), .Y(n227) );
  AO22X1_RVT U379 ( .A1(n666), .A2(\data_i[30][19] ), .A3(n665), .A4(
        \data_i[31][19] ), .Y(n226) );
  AO22X1_RVT U380 ( .A1(n668), .A2(\data_i[29][19] ), .A3(n667), .A4(
        \data_i[28][19] ), .Y(n225) );
  AO22X1_RVT U381 ( .A1(n674), .A2(\data_i[18][19] ), .A3(n673), .A4(
        \data_i[19][19] ), .Y(n232) );
  AO22X1_RVT U382 ( .A1(n676), .A2(\data_i[17][19] ), .A3(n675), .A4(
        \data_i[16][19] ), .Y(n231) );
  AO22X1_RVT U383 ( .A1(n678), .A2(\data_i[22][19] ), .A3(n677), .A4(
        \data_i[23][19] ), .Y(n230) );
  AO22X1_RVT U384 ( .A1(n680), .A2(\data_i[21][19] ), .A3(n679), .A4(
        \data_i[20][19] ), .Y(n229) );
  AO22X1_RVT U385 ( .A1(n638), .A2(\data_i[10][1] ), .A3(n637), .A4(
        \data_i[11][1] ), .Y(n240) );
  AO22X1_RVT U386 ( .A1(n640), .A2(\data_i[9][1] ), .A3(n639), .A4(
        \data_i[8][1] ), .Y(n239) );
  AO22X1_RVT U387 ( .A1(n642), .A2(\data_i[14][1] ), .A3(n641), .A4(
        \data_i[15][1] ), .Y(n238) );
  AO22X1_RVT U388 ( .A1(n644), .A2(\data_i[13][1] ), .A3(n643), .A4(
        \data_i[12][1] ), .Y(n237) );
  AO22X1_RVT U389 ( .A1(n650), .A2(\data_i[2][1] ), .A3(n649), .A4(
        \data_i[3][1] ), .Y(n244) );
  AO22X1_RVT U390 ( .A1(n652), .A2(\data_i[1][1] ), .A3(n651), .A4(
        \data_i[0][1] ), .Y(n243) );
  AO22X1_RVT U391 ( .A1(n654), .A2(\data_i[6][1] ), .A3(n653), .A4(
        \data_i[7][1] ), .Y(n242) );
  AO22X1_RVT U392 ( .A1(n656), .A2(\data_i[5][1] ), .A3(n655), .A4(
        \data_i[4][1] ), .Y(n241) );
  AO22X1_RVT U393 ( .A1(n662), .A2(\data_i[26][1] ), .A3(n661), .A4(
        \data_i[27][1] ), .Y(n248) );
  AO22X1_RVT U394 ( .A1(n664), .A2(\data_i[25][1] ), .A3(n663), .A4(
        \data_i[24][1] ), .Y(n247) );
  AO22X1_RVT U395 ( .A1(n666), .A2(\data_i[30][1] ), .A3(n665), .A4(
        \data_i[31][1] ), .Y(n246) );
  AO22X1_RVT U396 ( .A1(n668), .A2(\data_i[29][1] ), .A3(n667), .A4(
        \data_i[28][1] ), .Y(n245) );
  AO22X1_RVT U397 ( .A1(n674), .A2(\data_i[18][1] ), .A3(n673), .A4(
        \data_i[19][1] ), .Y(n252) );
  AO22X1_RVT U398 ( .A1(n676), .A2(\data_i[17][1] ), .A3(n675), .A4(
        \data_i[16][1] ), .Y(n251) );
  AO22X1_RVT U399 ( .A1(n678), .A2(\data_i[22][1] ), .A3(n677), .A4(
        \data_i[23][1] ), .Y(n250) );
  AO22X1_RVT U400 ( .A1(n680), .A2(\data_i[21][1] ), .A3(n679), .A4(
        \data_i[20][1] ), .Y(n249) );
  AO22X1_RVT U401 ( .A1(n638), .A2(\data_i[10][20] ), .A3(n637), .A4(
        \data_i[11][20] ), .Y(n260) );
  AO22X1_RVT U402 ( .A1(n640), .A2(\data_i[9][20] ), .A3(n639), .A4(
        \data_i[8][20] ), .Y(n259) );
  AO22X1_RVT U403 ( .A1(n642), .A2(\data_i[14][20] ), .A3(n641), .A4(
        \data_i[15][20] ), .Y(n258) );
  AO22X1_RVT U404 ( .A1(n644), .A2(\data_i[13][20] ), .A3(n643), .A4(
        \data_i[12][20] ), .Y(n257) );
  AO22X1_RVT U405 ( .A1(n650), .A2(\data_i[2][20] ), .A3(n649), .A4(
        \data_i[3][20] ), .Y(n264) );
  AO22X1_RVT U406 ( .A1(n652), .A2(\data_i[1][20] ), .A3(n651), .A4(
        \data_i[0][20] ), .Y(n263) );
  AO22X1_RVT U407 ( .A1(n654), .A2(\data_i[6][20] ), .A3(n653), .A4(
        \data_i[7][20] ), .Y(n262) );
  AO22X1_RVT U408 ( .A1(n656), .A2(\data_i[5][20] ), .A3(n655), .A4(
        \data_i[4][20] ), .Y(n261) );
  AO22X1_RVT U409 ( .A1(n662), .A2(\data_i[26][20] ), .A3(n661), .A4(
        \data_i[27][20] ), .Y(n268) );
  AO22X1_RVT U410 ( .A1(n664), .A2(\data_i[25][20] ), .A3(n663), .A4(
        \data_i[24][20] ), .Y(n267) );
  AO22X1_RVT U411 ( .A1(n666), .A2(\data_i[30][20] ), .A3(n665), .A4(
        \data_i[31][20] ), .Y(n266) );
  AO22X1_RVT U412 ( .A1(n668), .A2(\data_i[29][20] ), .A3(n667), .A4(
        \data_i[28][20] ), .Y(n265) );
  AO22X1_RVT U413 ( .A1(n674), .A2(\data_i[18][20] ), .A3(n673), .A4(
        \data_i[19][20] ), .Y(n272) );
  AO22X1_RVT U414 ( .A1(n676), .A2(\data_i[17][20] ), .A3(n675), .A4(
        \data_i[16][20] ), .Y(n271) );
  AO22X1_RVT U415 ( .A1(n678), .A2(\data_i[22][20] ), .A3(n677), .A4(
        \data_i[23][20] ), .Y(n270) );
  AO22X1_RVT U416 ( .A1(n680), .A2(\data_i[21][20] ), .A3(n679), .A4(
        \data_i[20][20] ), .Y(n269) );
  AO22X1_RVT U417 ( .A1(n638), .A2(\data_i[10][21] ), .A3(n637), .A4(
        \data_i[11][21] ), .Y(n280) );
  AO22X1_RVT U418 ( .A1(n640), .A2(\data_i[9][21] ), .A3(n639), .A4(
        \data_i[8][21] ), .Y(n279) );
  AO22X1_RVT U419 ( .A1(n642), .A2(\data_i[14][21] ), .A3(n641), .A4(
        \data_i[15][21] ), .Y(n278) );
  AO22X1_RVT U420 ( .A1(n644), .A2(\data_i[13][21] ), .A3(n643), .A4(
        \data_i[12][21] ), .Y(n277) );
  AO22X1_RVT U421 ( .A1(n650), .A2(\data_i[2][21] ), .A3(n649), .A4(
        \data_i[3][21] ), .Y(n284) );
  AO22X1_RVT U422 ( .A1(n652), .A2(\data_i[1][21] ), .A3(n651), .A4(
        \data_i[0][21] ), .Y(n283) );
  AO22X1_RVT U423 ( .A1(n654), .A2(\data_i[6][21] ), .A3(n653), .A4(
        \data_i[7][21] ), .Y(n282) );
  AO22X1_RVT U424 ( .A1(n656), .A2(\data_i[5][21] ), .A3(n655), .A4(
        \data_i[4][21] ), .Y(n281) );
  AO22X1_RVT U425 ( .A1(n662), .A2(\data_i[26][21] ), .A3(n661), .A4(
        \data_i[27][21] ), .Y(n288) );
  AO22X1_RVT U426 ( .A1(n664), .A2(\data_i[25][21] ), .A3(n663), .A4(
        \data_i[24][21] ), .Y(n287) );
  AO22X1_RVT U427 ( .A1(n666), .A2(\data_i[30][21] ), .A3(n665), .A4(
        \data_i[31][21] ), .Y(n286) );
  AO22X1_RVT U428 ( .A1(n668), .A2(\data_i[29][21] ), .A3(n667), .A4(
        \data_i[28][21] ), .Y(n285) );
  AO22X1_RVT U429 ( .A1(n674), .A2(\data_i[18][21] ), .A3(n673), .A4(
        \data_i[19][21] ), .Y(n292) );
  AO22X1_RVT U430 ( .A1(n676), .A2(\data_i[17][21] ), .A3(n675), .A4(
        \data_i[16][21] ), .Y(n291) );
  AO22X1_RVT U431 ( .A1(n678), .A2(\data_i[22][21] ), .A3(n677), .A4(
        \data_i[23][21] ), .Y(n290) );
  AO22X1_RVT U432 ( .A1(n680), .A2(\data_i[21][21] ), .A3(n679), .A4(
        \data_i[20][21] ), .Y(n289) );
  AO22X1_RVT U433 ( .A1(n638), .A2(\data_i[10][22] ), .A3(n637), .A4(
        \data_i[11][22] ), .Y(n300) );
  AO22X1_RVT U434 ( .A1(n640), .A2(\data_i[9][22] ), .A3(n639), .A4(
        \data_i[8][22] ), .Y(n299) );
  AO22X1_RVT U435 ( .A1(n642), .A2(\data_i[14][22] ), .A3(n641), .A4(
        \data_i[15][22] ), .Y(n298) );
  AO22X1_RVT U436 ( .A1(n644), .A2(\data_i[13][22] ), .A3(n643), .A4(
        \data_i[12][22] ), .Y(n297) );
  AO22X1_RVT U437 ( .A1(n650), .A2(\data_i[2][22] ), .A3(n649), .A4(
        \data_i[3][22] ), .Y(n304) );
  AO22X1_RVT U438 ( .A1(n652), .A2(\data_i[1][22] ), .A3(n651), .A4(
        \data_i[0][22] ), .Y(n303) );
  AO22X1_RVT U439 ( .A1(n654), .A2(\data_i[6][22] ), .A3(n653), .A4(
        \data_i[7][22] ), .Y(n302) );
  AO22X1_RVT U440 ( .A1(n656), .A2(\data_i[5][22] ), .A3(n655), .A4(
        \data_i[4][22] ), .Y(n301) );
  AO22X1_RVT U441 ( .A1(n662), .A2(\data_i[26][22] ), .A3(n661), .A4(
        \data_i[27][22] ), .Y(n308) );
  AO22X1_RVT U442 ( .A1(n664), .A2(\data_i[25][22] ), .A3(n663), .A4(
        \data_i[24][22] ), .Y(n307) );
  AO22X1_RVT U443 ( .A1(n666), .A2(\data_i[30][22] ), .A3(n665), .A4(
        \data_i[31][22] ), .Y(n306) );
  AO22X1_RVT U444 ( .A1(n668), .A2(\data_i[29][22] ), .A3(n667), .A4(
        \data_i[28][22] ), .Y(n305) );
  AO22X1_RVT U445 ( .A1(n674), .A2(\data_i[18][22] ), .A3(n673), .A4(
        \data_i[19][22] ), .Y(n312) );
  AO22X1_RVT U446 ( .A1(n676), .A2(\data_i[17][22] ), .A3(n675), .A4(
        \data_i[16][22] ), .Y(n311) );
  AO22X1_RVT U447 ( .A1(n678), .A2(\data_i[22][22] ), .A3(n677), .A4(
        \data_i[23][22] ), .Y(n310) );
  AO22X1_RVT U448 ( .A1(n680), .A2(\data_i[21][22] ), .A3(n679), .A4(
        \data_i[20][22] ), .Y(n309) );
  AO22X1_RVT U449 ( .A1(n638), .A2(\data_i[10][23] ), .A3(n637), .A4(
        \data_i[11][23] ), .Y(n320) );
  AO22X1_RVT U450 ( .A1(n640), .A2(\data_i[9][23] ), .A3(n639), .A4(
        \data_i[8][23] ), .Y(n319) );
  AO22X1_RVT U451 ( .A1(n642), .A2(\data_i[14][23] ), .A3(n641), .A4(
        \data_i[15][23] ), .Y(n318) );
  AO22X1_RVT U452 ( .A1(n644), .A2(\data_i[13][23] ), .A3(n643), .A4(
        \data_i[12][23] ), .Y(n317) );
  AO22X1_RVT U453 ( .A1(n650), .A2(\data_i[2][23] ), .A3(n649), .A4(
        \data_i[3][23] ), .Y(n324) );
  AO22X1_RVT U454 ( .A1(n652), .A2(\data_i[1][23] ), .A3(n651), .A4(
        \data_i[0][23] ), .Y(n323) );
  AO22X1_RVT U455 ( .A1(n654), .A2(\data_i[6][23] ), .A3(n653), .A4(
        \data_i[7][23] ), .Y(n322) );
  AO22X1_RVT U456 ( .A1(n656), .A2(\data_i[5][23] ), .A3(n655), .A4(
        \data_i[4][23] ), .Y(n321) );
  AO22X1_RVT U457 ( .A1(n662), .A2(\data_i[26][23] ), .A3(n661), .A4(
        \data_i[27][23] ), .Y(n328) );
  AO22X1_RVT U458 ( .A1(n664), .A2(\data_i[25][23] ), .A3(n663), .A4(
        \data_i[24][23] ), .Y(n327) );
  AO22X1_RVT U459 ( .A1(n666), .A2(\data_i[30][23] ), .A3(n665), .A4(
        \data_i[31][23] ), .Y(n326) );
  AO22X1_RVT U460 ( .A1(n668), .A2(\data_i[29][23] ), .A3(n667), .A4(
        \data_i[28][23] ), .Y(n325) );
  AO22X1_RVT U461 ( .A1(n674), .A2(\data_i[18][23] ), .A3(n673), .A4(
        \data_i[19][23] ), .Y(n332) );
  AO22X1_RVT U462 ( .A1(n676), .A2(\data_i[17][23] ), .A3(n675), .A4(
        \data_i[16][23] ), .Y(n331) );
  AO22X1_RVT U463 ( .A1(n678), .A2(\data_i[22][23] ), .A3(n677), .A4(
        \data_i[23][23] ), .Y(n330) );
  AO22X1_RVT U464 ( .A1(n680), .A2(\data_i[21][23] ), .A3(n679), .A4(
        \data_i[20][23] ), .Y(n329) );
  AO22X1_RVT U465 ( .A1(n638), .A2(\data_i[10][24] ), .A3(n637), .A4(
        \data_i[11][24] ), .Y(n340) );
  AO22X1_RVT U466 ( .A1(n640), .A2(\data_i[9][24] ), .A3(n639), .A4(
        \data_i[8][24] ), .Y(n339) );
  AO22X1_RVT U467 ( .A1(n642), .A2(\data_i[14][24] ), .A3(n641), .A4(
        \data_i[15][24] ), .Y(n338) );
  AO22X1_RVT U468 ( .A1(n644), .A2(\data_i[13][24] ), .A3(n643), .A4(
        \data_i[12][24] ), .Y(n337) );
  AO22X1_RVT U469 ( .A1(n650), .A2(\data_i[2][24] ), .A3(n649), .A4(
        \data_i[3][24] ), .Y(n344) );
  AO22X1_RVT U470 ( .A1(n652), .A2(\data_i[1][24] ), .A3(n651), .A4(
        \data_i[0][24] ), .Y(n343) );
  AO22X1_RVT U471 ( .A1(n654), .A2(\data_i[6][24] ), .A3(n653), .A4(
        \data_i[7][24] ), .Y(n342) );
  AO22X1_RVT U472 ( .A1(n656), .A2(\data_i[5][24] ), .A3(n655), .A4(
        \data_i[4][24] ), .Y(n341) );
  AO22X1_RVT U473 ( .A1(n662), .A2(\data_i[26][24] ), .A3(n661), .A4(
        \data_i[27][24] ), .Y(n348) );
  AO22X1_RVT U474 ( .A1(n664), .A2(\data_i[25][24] ), .A3(n663), .A4(
        \data_i[24][24] ), .Y(n347) );
  AO22X1_RVT U475 ( .A1(n666), .A2(\data_i[30][24] ), .A3(n665), .A4(
        \data_i[31][24] ), .Y(n346) );
  AO22X1_RVT U476 ( .A1(n668), .A2(\data_i[29][24] ), .A3(n667), .A4(
        \data_i[28][24] ), .Y(n345) );
  AO22X1_RVT U477 ( .A1(n674), .A2(\data_i[18][24] ), .A3(n673), .A4(
        \data_i[19][24] ), .Y(n352) );
  AO22X1_RVT U478 ( .A1(n676), .A2(\data_i[17][24] ), .A3(n675), .A4(
        \data_i[16][24] ), .Y(n351) );
  AO22X1_RVT U479 ( .A1(n678), .A2(\data_i[22][24] ), .A3(n677), .A4(
        \data_i[23][24] ), .Y(n350) );
  AO22X1_RVT U480 ( .A1(n680), .A2(\data_i[21][24] ), .A3(n679), .A4(
        \data_i[20][24] ), .Y(n349) );
  AO22X1_RVT U481 ( .A1(n638), .A2(\data_i[10][25] ), .A3(n637), .A4(
        \data_i[11][25] ), .Y(n360) );
  AO22X1_RVT U482 ( .A1(n640), .A2(\data_i[9][25] ), .A3(n639), .A4(
        \data_i[8][25] ), .Y(n359) );
  AO22X1_RVT U483 ( .A1(n642), .A2(\data_i[14][25] ), .A3(n641), .A4(
        \data_i[15][25] ), .Y(n358) );
  AO22X1_RVT U484 ( .A1(n644), .A2(\data_i[13][25] ), .A3(n643), .A4(
        \data_i[12][25] ), .Y(n357) );
  AO22X1_RVT U485 ( .A1(n650), .A2(\data_i[2][25] ), .A3(n649), .A4(
        \data_i[3][25] ), .Y(n364) );
  AO22X1_RVT U486 ( .A1(n652), .A2(\data_i[1][25] ), .A3(n651), .A4(
        \data_i[0][25] ), .Y(n363) );
  AO22X1_RVT U487 ( .A1(n654), .A2(\data_i[6][25] ), .A3(n653), .A4(
        \data_i[7][25] ), .Y(n362) );
  AO22X1_RVT U488 ( .A1(n656), .A2(\data_i[5][25] ), .A3(n655), .A4(
        \data_i[4][25] ), .Y(n361) );
  AO22X1_RVT U489 ( .A1(n662), .A2(\data_i[26][25] ), .A3(n661), .A4(
        \data_i[27][25] ), .Y(n368) );
  AO22X1_RVT U490 ( .A1(n664), .A2(\data_i[25][25] ), .A3(n663), .A4(
        \data_i[24][25] ), .Y(n367) );
  AO22X1_RVT U491 ( .A1(n666), .A2(\data_i[30][25] ), .A3(n665), .A4(
        \data_i[31][25] ), .Y(n366) );
  AO22X1_RVT U492 ( .A1(n668), .A2(\data_i[29][25] ), .A3(n667), .A4(
        \data_i[28][25] ), .Y(n365) );
  AO22X1_RVT U493 ( .A1(n674), .A2(\data_i[18][25] ), .A3(n673), .A4(
        \data_i[19][25] ), .Y(n372) );
  AO22X1_RVT U494 ( .A1(n676), .A2(\data_i[17][25] ), .A3(n675), .A4(
        \data_i[16][25] ), .Y(n371) );
  AO22X1_RVT U495 ( .A1(n678), .A2(\data_i[22][25] ), .A3(n677), .A4(
        \data_i[23][25] ), .Y(n370) );
  AO22X1_RVT U496 ( .A1(n680), .A2(\data_i[21][25] ), .A3(n679), .A4(
        \data_i[20][25] ), .Y(n369) );
  AO22X1_RVT U497 ( .A1(n638), .A2(\data_i[10][26] ), .A3(n637), .A4(
        \data_i[11][26] ), .Y(n380) );
  AO22X1_RVT U498 ( .A1(n640), .A2(\data_i[9][26] ), .A3(n639), .A4(
        \data_i[8][26] ), .Y(n379) );
  AO22X1_RVT U499 ( .A1(n642), .A2(\data_i[14][26] ), .A3(n641), .A4(
        \data_i[15][26] ), .Y(n378) );
  AO22X1_RVT U500 ( .A1(n644), .A2(\data_i[13][26] ), .A3(n643), .A4(
        \data_i[12][26] ), .Y(n377) );
  AO22X1_RVT U501 ( .A1(n650), .A2(\data_i[2][26] ), .A3(n649), .A4(
        \data_i[3][26] ), .Y(n384) );
  AO22X1_RVT U502 ( .A1(n652), .A2(\data_i[1][26] ), .A3(n651), .A4(
        \data_i[0][26] ), .Y(n383) );
  AO22X1_RVT U503 ( .A1(n654), .A2(\data_i[6][26] ), .A3(n653), .A4(
        \data_i[7][26] ), .Y(n382) );
  AO22X1_RVT U504 ( .A1(n656), .A2(\data_i[5][26] ), .A3(n655), .A4(
        \data_i[4][26] ), .Y(n381) );
  AO22X1_RVT U505 ( .A1(n662), .A2(\data_i[26][26] ), .A3(n661), .A4(
        \data_i[27][26] ), .Y(n388) );
  AO22X1_RVT U506 ( .A1(n664), .A2(\data_i[25][26] ), .A3(n663), .A4(
        \data_i[24][26] ), .Y(n387) );
  AO22X1_RVT U507 ( .A1(n666), .A2(\data_i[30][26] ), .A3(n665), .A4(
        \data_i[31][26] ), .Y(n386) );
  AO22X1_RVT U508 ( .A1(n668), .A2(\data_i[29][26] ), .A3(n667), .A4(
        \data_i[28][26] ), .Y(n385) );
  AO22X1_RVT U509 ( .A1(n674), .A2(\data_i[18][26] ), .A3(n673), .A4(
        \data_i[19][26] ), .Y(n392) );
  AO22X1_RVT U510 ( .A1(n676), .A2(\data_i[17][26] ), .A3(n675), .A4(
        \data_i[16][26] ), .Y(n391) );
  AO22X1_RVT U511 ( .A1(n678), .A2(\data_i[22][26] ), .A3(n677), .A4(
        \data_i[23][26] ), .Y(n390) );
  AO22X1_RVT U512 ( .A1(n680), .A2(\data_i[21][26] ), .A3(n679), .A4(
        \data_i[20][26] ), .Y(n389) );
  AO22X1_RVT U513 ( .A1(n638), .A2(\data_i[10][27] ), .A3(n637), .A4(
        \data_i[11][27] ), .Y(n400) );
  AO22X1_RVT U514 ( .A1(n640), .A2(\data_i[9][27] ), .A3(n639), .A4(
        \data_i[8][27] ), .Y(n399) );
  AO22X1_RVT U515 ( .A1(n642), .A2(\data_i[14][27] ), .A3(n641), .A4(
        \data_i[15][27] ), .Y(n398) );
  AO22X1_RVT U516 ( .A1(n644), .A2(\data_i[13][27] ), .A3(n643), .A4(
        \data_i[12][27] ), .Y(n397) );
  AO22X1_RVT U517 ( .A1(n650), .A2(\data_i[2][27] ), .A3(n649), .A4(
        \data_i[3][27] ), .Y(n404) );
  AO22X1_RVT U518 ( .A1(n652), .A2(\data_i[1][27] ), .A3(n651), .A4(
        \data_i[0][27] ), .Y(n403) );
  AO22X1_RVT U519 ( .A1(n654), .A2(\data_i[6][27] ), .A3(n653), .A4(
        \data_i[7][27] ), .Y(n402) );
  AO22X1_RVT U520 ( .A1(n656), .A2(\data_i[5][27] ), .A3(n655), .A4(
        \data_i[4][27] ), .Y(n401) );
  AO22X1_RVT U521 ( .A1(n662), .A2(\data_i[26][27] ), .A3(n661), .A4(
        \data_i[27][27] ), .Y(n408) );
  AO22X1_RVT U522 ( .A1(n664), .A2(\data_i[25][27] ), .A3(n663), .A4(
        \data_i[24][27] ), .Y(n407) );
  AO22X1_RVT U523 ( .A1(n666), .A2(\data_i[30][27] ), .A3(n665), .A4(
        \data_i[31][27] ), .Y(n406) );
  AO22X1_RVT U524 ( .A1(n668), .A2(\data_i[29][27] ), .A3(n667), .A4(
        \data_i[28][27] ), .Y(n405) );
  AO22X1_RVT U525 ( .A1(n674), .A2(\data_i[18][27] ), .A3(n673), .A4(
        \data_i[19][27] ), .Y(n412) );
  AO22X1_RVT U526 ( .A1(n676), .A2(\data_i[17][27] ), .A3(n675), .A4(
        \data_i[16][27] ), .Y(n411) );
  AO22X1_RVT U527 ( .A1(n678), .A2(\data_i[22][27] ), .A3(n677), .A4(
        \data_i[23][27] ), .Y(n410) );
  AO22X1_RVT U528 ( .A1(n680), .A2(\data_i[21][27] ), .A3(n679), .A4(
        \data_i[20][27] ), .Y(n409) );
  AO22X1_RVT U529 ( .A1(n638), .A2(\data_i[10][28] ), .A3(n637), .A4(
        \data_i[11][28] ), .Y(n420) );
  AO22X1_RVT U530 ( .A1(n640), .A2(\data_i[9][28] ), .A3(n639), .A4(
        \data_i[8][28] ), .Y(n419) );
  AO22X1_RVT U531 ( .A1(n642), .A2(\data_i[14][28] ), .A3(n641), .A4(
        \data_i[15][28] ), .Y(n418) );
  AO22X1_RVT U532 ( .A1(n644), .A2(\data_i[13][28] ), .A3(n643), .A4(
        \data_i[12][28] ), .Y(n417) );
  AO22X1_RVT U533 ( .A1(n650), .A2(\data_i[2][28] ), .A3(n649), .A4(
        \data_i[3][28] ), .Y(n424) );
  AO22X1_RVT U534 ( .A1(n652), .A2(\data_i[1][28] ), .A3(n651), .A4(
        \data_i[0][28] ), .Y(n423) );
  AO22X1_RVT U535 ( .A1(n654), .A2(\data_i[6][28] ), .A3(n653), .A4(
        \data_i[7][28] ), .Y(n422) );
  AO22X1_RVT U536 ( .A1(n656), .A2(\data_i[5][28] ), .A3(n655), .A4(
        \data_i[4][28] ), .Y(n421) );
  AO22X1_RVT U537 ( .A1(n662), .A2(\data_i[26][28] ), .A3(n661), .A4(
        \data_i[27][28] ), .Y(n428) );
  AO22X1_RVT U538 ( .A1(n664), .A2(\data_i[25][28] ), .A3(n663), .A4(
        \data_i[24][28] ), .Y(n427) );
  AO22X1_RVT U539 ( .A1(n666), .A2(\data_i[30][28] ), .A3(n665), .A4(
        \data_i[31][28] ), .Y(n426) );
  AO22X1_RVT U540 ( .A1(n668), .A2(\data_i[29][28] ), .A3(n667), .A4(
        \data_i[28][28] ), .Y(n425) );
  AO22X1_RVT U541 ( .A1(n674), .A2(\data_i[18][28] ), .A3(n673), .A4(
        \data_i[19][28] ), .Y(n432) );
  AO22X1_RVT U542 ( .A1(n676), .A2(\data_i[17][28] ), .A3(n675), .A4(
        \data_i[16][28] ), .Y(n431) );
  AO22X1_RVT U543 ( .A1(n678), .A2(\data_i[22][28] ), .A3(n677), .A4(
        \data_i[23][28] ), .Y(n430) );
  AO22X1_RVT U544 ( .A1(n680), .A2(\data_i[21][28] ), .A3(n679), .A4(
        \data_i[20][28] ), .Y(n429) );
  AO22X1_RVT U545 ( .A1(n638), .A2(\data_i[10][29] ), .A3(n637), .A4(
        \data_i[11][29] ), .Y(n440) );
  AO22X1_RVT U546 ( .A1(n640), .A2(\data_i[9][29] ), .A3(n639), .A4(
        \data_i[8][29] ), .Y(n439) );
  AO22X1_RVT U547 ( .A1(n642), .A2(\data_i[14][29] ), .A3(n641), .A4(
        \data_i[15][29] ), .Y(n438) );
  AO22X1_RVT U548 ( .A1(n644), .A2(\data_i[13][29] ), .A3(n643), .A4(
        \data_i[12][29] ), .Y(n437) );
  AO22X1_RVT U549 ( .A1(n650), .A2(\data_i[2][29] ), .A3(n649), .A4(
        \data_i[3][29] ), .Y(n444) );
  AO22X1_RVT U550 ( .A1(n652), .A2(\data_i[1][29] ), .A3(n651), .A4(
        \data_i[0][29] ), .Y(n443) );
  AO22X1_RVT U551 ( .A1(n654), .A2(\data_i[6][29] ), .A3(n653), .A4(
        \data_i[7][29] ), .Y(n442) );
  AO22X1_RVT U552 ( .A1(n656), .A2(\data_i[5][29] ), .A3(n655), .A4(
        \data_i[4][29] ), .Y(n441) );
  AO22X1_RVT U553 ( .A1(n662), .A2(\data_i[26][29] ), .A3(n661), .A4(
        \data_i[27][29] ), .Y(n448) );
  AO22X1_RVT U554 ( .A1(n664), .A2(\data_i[25][29] ), .A3(n663), .A4(
        \data_i[24][29] ), .Y(n447) );
  AO22X1_RVT U555 ( .A1(n666), .A2(\data_i[30][29] ), .A3(n665), .A4(
        \data_i[31][29] ), .Y(n446) );
  AO22X1_RVT U556 ( .A1(n668), .A2(\data_i[29][29] ), .A3(n667), .A4(
        \data_i[28][29] ), .Y(n445) );
  AO22X1_RVT U557 ( .A1(n674), .A2(\data_i[18][29] ), .A3(n673), .A4(
        \data_i[19][29] ), .Y(n452) );
  AO22X1_RVT U558 ( .A1(n676), .A2(\data_i[17][29] ), .A3(n675), .A4(
        \data_i[16][29] ), .Y(n451) );
  AO22X1_RVT U559 ( .A1(n678), .A2(\data_i[22][29] ), .A3(n677), .A4(
        \data_i[23][29] ), .Y(n450) );
  AO22X1_RVT U560 ( .A1(n680), .A2(\data_i[21][29] ), .A3(n679), .A4(
        \data_i[20][29] ), .Y(n449) );
  AO22X1_RVT U561 ( .A1(n638), .A2(\data_i[10][2] ), .A3(n637), .A4(
        \data_i[11][2] ), .Y(n460) );
  AO22X1_RVT U562 ( .A1(n640), .A2(\data_i[9][2] ), .A3(n639), .A4(
        \data_i[8][2] ), .Y(n459) );
  AO22X1_RVT U563 ( .A1(n642), .A2(\data_i[14][2] ), .A3(n641), .A4(
        \data_i[15][2] ), .Y(n458) );
  AO22X1_RVT U564 ( .A1(n644), .A2(\data_i[13][2] ), .A3(n643), .A4(
        \data_i[12][2] ), .Y(n457) );
  AO22X1_RVT U565 ( .A1(n650), .A2(\data_i[2][2] ), .A3(n649), .A4(
        \data_i[3][2] ), .Y(n464) );
  AO22X1_RVT U566 ( .A1(n652), .A2(\data_i[1][2] ), .A3(n651), .A4(
        \data_i[0][2] ), .Y(n463) );
  AO22X1_RVT U567 ( .A1(n654), .A2(\data_i[6][2] ), .A3(n653), .A4(
        \data_i[7][2] ), .Y(n462) );
  AO22X1_RVT U568 ( .A1(n656), .A2(\data_i[5][2] ), .A3(n655), .A4(
        \data_i[4][2] ), .Y(n461) );
  AO22X1_RVT U569 ( .A1(n662), .A2(\data_i[26][2] ), .A3(n661), .A4(
        \data_i[27][2] ), .Y(n468) );
  AO22X1_RVT U570 ( .A1(n664), .A2(\data_i[25][2] ), .A3(n663), .A4(
        \data_i[24][2] ), .Y(n467) );
  AO22X1_RVT U571 ( .A1(n666), .A2(\data_i[30][2] ), .A3(n665), .A4(
        \data_i[31][2] ), .Y(n466) );
  AO22X1_RVT U572 ( .A1(n668), .A2(\data_i[29][2] ), .A3(n667), .A4(
        \data_i[28][2] ), .Y(n465) );
  AO22X1_RVT U573 ( .A1(n674), .A2(\data_i[18][2] ), .A3(n673), .A4(
        \data_i[19][2] ), .Y(n472) );
  AO22X1_RVT U574 ( .A1(n676), .A2(\data_i[17][2] ), .A3(n675), .A4(
        \data_i[16][2] ), .Y(n471) );
  AO22X1_RVT U575 ( .A1(n678), .A2(\data_i[22][2] ), .A3(n677), .A4(
        \data_i[23][2] ), .Y(n470) );
  AO22X1_RVT U576 ( .A1(n680), .A2(\data_i[21][2] ), .A3(n679), .A4(
        \data_i[20][2] ), .Y(n469) );
  AO22X1_RVT U577 ( .A1(n638), .A2(\data_i[10][30] ), .A3(n637), .A4(
        \data_i[11][30] ), .Y(n480) );
  AO22X1_RVT U578 ( .A1(n640), .A2(\data_i[9][30] ), .A3(n639), .A4(
        \data_i[8][30] ), .Y(n479) );
  AO22X1_RVT U579 ( .A1(n642), .A2(\data_i[14][30] ), .A3(n641), .A4(
        \data_i[15][30] ), .Y(n478) );
  AO22X1_RVT U580 ( .A1(n644), .A2(\data_i[13][30] ), .A3(n643), .A4(
        \data_i[12][30] ), .Y(n477) );
  AO22X1_RVT U581 ( .A1(n650), .A2(\data_i[2][30] ), .A3(n649), .A4(
        \data_i[3][30] ), .Y(n484) );
  AO22X1_RVT U582 ( .A1(n652), .A2(\data_i[1][30] ), .A3(n651), .A4(
        \data_i[0][30] ), .Y(n483) );
  AO22X1_RVT U583 ( .A1(n654), .A2(\data_i[6][30] ), .A3(n653), .A4(
        \data_i[7][30] ), .Y(n482) );
  AO22X1_RVT U584 ( .A1(n656), .A2(\data_i[5][30] ), .A3(n655), .A4(
        \data_i[4][30] ), .Y(n481) );
  AO22X1_RVT U585 ( .A1(n662), .A2(\data_i[26][30] ), .A3(n661), .A4(
        \data_i[27][30] ), .Y(n488) );
  AO22X1_RVT U586 ( .A1(n664), .A2(\data_i[25][30] ), .A3(n663), .A4(
        \data_i[24][30] ), .Y(n487) );
  AO22X1_RVT U587 ( .A1(n666), .A2(\data_i[30][30] ), .A3(n665), .A4(
        \data_i[31][30] ), .Y(n486) );
  AO22X1_RVT U588 ( .A1(n668), .A2(\data_i[29][30] ), .A3(n667), .A4(
        \data_i[28][30] ), .Y(n485) );
  AO22X1_RVT U589 ( .A1(n674), .A2(\data_i[18][30] ), .A3(n673), .A4(
        \data_i[19][30] ), .Y(n492) );
  AO22X1_RVT U590 ( .A1(n676), .A2(\data_i[17][30] ), .A3(n675), .A4(
        \data_i[16][30] ), .Y(n491) );
  AO22X1_RVT U591 ( .A1(n678), .A2(\data_i[22][30] ), .A3(n677), .A4(
        \data_i[23][30] ), .Y(n490) );
  AO22X1_RVT U592 ( .A1(n680), .A2(\data_i[21][30] ), .A3(n679), .A4(
        \data_i[20][30] ), .Y(n489) );
  AO22X1_RVT U593 ( .A1(n638), .A2(\data_i[10][31] ), .A3(n637), .A4(
        \data_i[11][31] ), .Y(n500) );
  AO22X1_RVT U594 ( .A1(n640), .A2(\data_i[9][31] ), .A3(n639), .A4(
        \data_i[8][31] ), .Y(n499) );
  AO22X1_RVT U595 ( .A1(n642), .A2(\data_i[14][31] ), .A3(n641), .A4(
        \data_i[15][31] ), .Y(n498) );
  AO22X1_RVT U596 ( .A1(n644), .A2(\data_i[13][31] ), .A3(n643), .A4(
        \data_i[12][31] ), .Y(n497) );
  AO22X1_RVT U597 ( .A1(n650), .A2(\data_i[2][31] ), .A3(n649), .A4(
        \data_i[3][31] ), .Y(n504) );
  AO22X1_RVT U598 ( .A1(n652), .A2(\data_i[1][31] ), .A3(n651), .A4(
        \data_i[0][31] ), .Y(n503) );
  AO22X1_RVT U599 ( .A1(n654), .A2(\data_i[6][31] ), .A3(n653), .A4(
        \data_i[7][31] ), .Y(n502) );
  AO22X1_RVT U600 ( .A1(n656), .A2(\data_i[5][31] ), .A3(n655), .A4(
        \data_i[4][31] ), .Y(n501) );
  AO22X1_RVT U601 ( .A1(n662), .A2(\data_i[26][31] ), .A3(n661), .A4(
        \data_i[27][31] ), .Y(n508) );
  AO22X1_RVT U602 ( .A1(n664), .A2(\data_i[25][31] ), .A3(n663), .A4(
        \data_i[24][31] ), .Y(n507) );
  AO22X1_RVT U603 ( .A1(n666), .A2(\data_i[30][31] ), .A3(n665), .A4(
        \data_i[31][31] ), .Y(n506) );
  AO22X1_RVT U604 ( .A1(n668), .A2(\data_i[29][31] ), .A3(n667), .A4(
        \data_i[28][31] ), .Y(n505) );
  AO22X1_RVT U605 ( .A1(n674), .A2(\data_i[18][31] ), .A3(n673), .A4(
        \data_i[19][31] ), .Y(n512) );
  AO22X1_RVT U606 ( .A1(n676), .A2(\data_i[17][31] ), .A3(n675), .A4(
        \data_i[16][31] ), .Y(n511) );
  AO22X1_RVT U607 ( .A1(n678), .A2(\data_i[22][31] ), .A3(n677), .A4(
        \data_i[23][31] ), .Y(n510) );
  AO22X1_RVT U608 ( .A1(n680), .A2(\data_i[21][31] ), .A3(n679), .A4(
        \data_i[20][31] ), .Y(n509) );
  AO22X1_RVT U609 ( .A1(n638), .A2(\data_i[10][3] ), .A3(n637), .A4(
        \data_i[11][3] ), .Y(n520) );
  AO22X1_RVT U610 ( .A1(n640), .A2(\data_i[9][3] ), .A3(n639), .A4(
        \data_i[8][3] ), .Y(n519) );
  AO22X1_RVT U611 ( .A1(n642), .A2(\data_i[14][3] ), .A3(n641), .A4(
        \data_i[15][3] ), .Y(n518) );
  AO22X1_RVT U612 ( .A1(n644), .A2(\data_i[13][3] ), .A3(n643), .A4(
        \data_i[12][3] ), .Y(n517) );
  AO22X1_RVT U613 ( .A1(n650), .A2(\data_i[2][3] ), .A3(n649), .A4(
        \data_i[3][3] ), .Y(n524) );
  AO22X1_RVT U614 ( .A1(n652), .A2(\data_i[1][3] ), .A3(n651), .A4(
        \data_i[0][3] ), .Y(n523) );
  AO22X1_RVT U615 ( .A1(n654), .A2(\data_i[6][3] ), .A3(n653), .A4(
        \data_i[7][3] ), .Y(n522) );
  AO22X1_RVT U616 ( .A1(n656), .A2(\data_i[5][3] ), .A3(n655), .A4(
        \data_i[4][3] ), .Y(n521) );
  AO22X1_RVT U617 ( .A1(n662), .A2(\data_i[26][3] ), .A3(n661), .A4(
        \data_i[27][3] ), .Y(n528) );
  AO22X1_RVT U618 ( .A1(n664), .A2(\data_i[25][3] ), .A3(n663), .A4(
        \data_i[24][3] ), .Y(n527) );
  AO22X1_RVT U619 ( .A1(n666), .A2(\data_i[30][3] ), .A3(n665), .A4(
        \data_i[31][3] ), .Y(n526) );
  AO22X1_RVT U620 ( .A1(n668), .A2(\data_i[29][3] ), .A3(n667), .A4(
        \data_i[28][3] ), .Y(n525) );
  AO22X1_RVT U621 ( .A1(n674), .A2(\data_i[18][3] ), .A3(n673), .A4(
        \data_i[19][3] ), .Y(n532) );
  AO22X1_RVT U622 ( .A1(n676), .A2(\data_i[17][3] ), .A3(n675), .A4(
        \data_i[16][3] ), .Y(n531) );
  AO22X1_RVT U623 ( .A1(n678), .A2(\data_i[22][3] ), .A3(n677), .A4(
        \data_i[23][3] ), .Y(n530) );
  AO22X1_RVT U624 ( .A1(n680), .A2(\data_i[21][3] ), .A3(n679), .A4(
        \data_i[20][3] ), .Y(n529) );
  AO22X1_RVT U625 ( .A1(n638), .A2(\data_i[10][4] ), .A3(n637), .A4(
        \data_i[11][4] ), .Y(n540) );
  AO22X1_RVT U626 ( .A1(n640), .A2(\data_i[9][4] ), .A3(n639), .A4(
        \data_i[8][4] ), .Y(n539) );
  AO22X1_RVT U627 ( .A1(n642), .A2(\data_i[14][4] ), .A3(n641), .A4(
        \data_i[15][4] ), .Y(n538) );
  AO22X1_RVT U628 ( .A1(n644), .A2(\data_i[13][4] ), .A3(n643), .A4(
        \data_i[12][4] ), .Y(n537) );
  AO22X1_RVT U629 ( .A1(n650), .A2(\data_i[2][4] ), .A3(n649), .A4(
        \data_i[3][4] ), .Y(n544) );
  AO22X1_RVT U630 ( .A1(n652), .A2(\data_i[1][4] ), .A3(n651), .A4(
        \data_i[0][4] ), .Y(n543) );
  AO22X1_RVT U631 ( .A1(n654), .A2(\data_i[6][4] ), .A3(n653), .A4(
        \data_i[7][4] ), .Y(n542) );
  AO22X1_RVT U632 ( .A1(n656), .A2(\data_i[5][4] ), .A3(n655), .A4(
        \data_i[4][4] ), .Y(n541) );
  AO22X1_RVT U633 ( .A1(n662), .A2(\data_i[26][4] ), .A3(n661), .A4(
        \data_i[27][4] ), .Y(n548) );
  AO22X1_RVT U634 ( .A1(n664), .A2(\data_i[25][4] ), .A3(n663), .A4(
        \data_i[24][4] ), .Y(n547) );
  AO22X1_RVT U635 ( .A1(n666), .A2(\data_i[30][4] ), .A3(n665), .A4(
        \data_i[31][4] ), .Y(n546) );
  AO22X1_RVT U636 ( .A1(n668), .A2(\data_i[29][4] ), .A3(n667), .A4(
        \data_i[28][4] ), .Y(n545) );
  AO22X1_RVT U637 ( .A1(n674), .A2(\data_i[18][4] ), .A3(n673), .A4(
        \data_i[19][4] ), .Y(n552) );
  AO22X1_RVT U638 ( .A1(n676), .A2(\data_i[17][4] ), .A3(n675), .A4(
        \data_i[16][4] ), .Y(n551) );
  AO22X1_RVT U639 ( .A1(n678), .A2(\data_i[22][4] ), .A3(n677), .A4(
        \data_i[23][4] ), .Y(n550) );
  AO22X1_RVT U640 ( .A1(n680), .A2(\data_i[21][4] ), .A3(n679), .A4(
        \data_i[20][4] ), .Y(n549) );
  AO22X1_RVT U641 ( .A1(n638), .A2(\data_i[10][5] ), .A3(n637), .A4(
        \data_i[11][5] ), .Y(n560) );
  AO22X1_RVT U642 ( .A1(n640), .A2(\data_i[9][5] ), .A3(n639), .A4(
        \data_i[8][5] ), .Y(n559) );
  AO22X1_RVT U643 ( .A1(n642), .A2(\data_i[14][5] ), .A3(n641), .A4(
        \data_i[15][5] ), .Y(n558) );
  AO22X1_RVT U644 ( .A1(n644), .A2(\data_i[13][5] ), .A3(n643), .A4(
        \data_i[12][5] ), .Y(n557) );
  AO22X1_RVT U645 ( .A1(n650), .A2(\data_i[2][5] ), .A3(n649), .A4(
        \data_i[3][5] ), .Y(n564) );
  AO22X1_RVT U646 ( .A1(n652), .A2(\data_i[1][5] ), .A3(n651), .A4(
        \data_i[0][5] ), .Y(n563) );
  AO22X1_RVT U647 ( .A1(n654), .A2(\data_i[6][5] ), .A3(n653), .A4(
        \data_i[7][5] ), .Y(n562) );
  AO22X1_RVT U648 ( .A1(n656), .A2(\data_i[5][5] ), .A3(n655), .A4(
        \data_i[4][5] ), .Y(n561) );
  AO22X1_RVT U649 ( .A1(n662), .A2(\data_i[26][5] ), .A3(n661), .A4(
        \data_i[27][5] ), .Y(n568) );
  AO22X1_RVT U650 ( .A1(n664), .A2(\data_i[25][5] ), .A3(n663), .A4(
        \data_i[24][5] ), .Y(n567) );
  AO22X1_RVT U651 ( .A1(n666), .A2(\data_i[30][5] ), .A3(n665), .A4(
        \data_i[31][5] ), .Y(n566) );
  AO22X1_RVT U652 ( .A1(n668), .A2(\data_i[29][5] ), .A3(n667), .A4(
        \data_i[28][5] ), .Y(n565) );
  AO22X1_RVT U653 ( .A1(n674), .A2(\data_i[18][5] ), .A3(n673), .A4(
        \data_i[19][5] ), .Y(n572) );
  AO22X1_RVT U654 ( .A1(n676), .A2(\data_i[17][5] ), .A3(n675), .A4(
        \data_i[16][5] ), .Y(n571) );
  AO22X1_RVT U655 ( .A1(n678), .A2(\data_i[22][5] ), .A3(n677), .A4(
        \data_i[23][5] ), .Y(n570) );
  AO22X1_RVT U656 ( .A1(n680), .A2(\data_i[21][5] ), .A3(n679), .A4(
        \data_i[20][5] ), .Y(n569) );
  AO22X1_RVT U657 ( .A1(n638), .A2(\data_i[10][6] ), .A3(n637), .A4(
        \data_i[11][6] ), .Y(n580) );
  AO22X1_RVT U658 ( .A1(n640), .A2(\data_i[9][6] ), .A3(n639), .A4(
        \data_i[8][6] ), .Y(n579) );
  AO22X1_RVT U659 ( .A1(n642), .A2(\data_i[14][6] ), .A3(n641), .A4(
        \data_i[15][6] ), .Y(n578) );
  AO22X1_RVT U660 ( .A1(n644), .A2(\data_i[13][6] ), .A3(n643), .A4(
        \data_i[12][6] ), .Y(n577) );
  AO22X1_RVT U661 ( .A1(n650), .A2(\data_i[2][6] ), .A3(n649), .A4(
        \data_i[3][6] ), .Y(n584) );
  AO22X1_RVT U662 ( .A1(n652), .A2(\data_i[1][6] ), .A3(n651), .A4(
        \data_i[0][6] ), .Y(n583) );
  AO22X1_RVT U663 ( .A1(n654), .A2(\data_i[6][6] ), .A3(n653), .A4(
        \data_i[7][6] ), .Y(n582) );
  AO22X1_RVT U664 ( .A1(n656), .A2(\data_i[5][6] ), .A3(n655), .A4(
        \data_i[4][6] ), .Y(n581) );
  AO22X1_RVT U665 ( .A1(n662), .A2(\data_i[26][6] ), .A3(n661), .A4(
        \data_i[27][6] ), .Y(n588) );
  AO22X1_RVT U666 ( .A1(n664), .A2(\data_i[25][6] ), .A3(n663), .A4(
        \data_i[24][6] ), .Y(n587) );
  AO22X1_RVT U667 ( .A1(n666), .A2(\data_i[30][6] ), .A3(n665), .A4(
        \data_i[31][6] ), .Y(n586) );
  AO22X1_RVT U668 ( .A1(n668), .A2(\data_i[29][6] ), .A3(n667), .A4(
        \data_i[28][6] ), .Y(n585) );
  AO22X1_RVT U669 ( .A1(n674), .A2(\data_i[18][6] ), .A3(n673), .A4(
        \data_i[19][6] ), .Y(n592) );
  AO22X1_RVT U670 ( .A1(n676), .A2(\data_i[17][6] ), .A3(n675), .A4(
        \data_i[16][6] ), .Y(n591) );
  AO22X1_RVT U671 ( .A1(n678), .A2(\data_i[22][6] ), .A3(n677), .A4(
        \data_i[23][6] ), .Y(n590) );
  AO22X1_RVT U672 ( .A1(n680), .A2(\data_i[21][6] ), .A3(n679), .A4(
        \data_i[20][6] ), .Y(n589) );
  AO22X1_RVT U673 ( .A1(n638), .A2(\data_i[10][7] ), .A3(n637), .A4(
        \data_i[11][7] ), .Y(n600) );
  AO22X1_RVT U674 ( .A1(n640), .A2(\data_i[9][7] ), .A3(n639), .A4(
        \data_i[8][7] ), .Y(n599) );
  AO22X1_RVT U675 ( .A1(n642), .A2(\data_i[14][7] ), .A3(n641), .A4(
        \data_i[15][7] ), .Y(n598) );
  AO22X1_RVT U676 ( .A1(n644), .A2(\data_i[13][7] ), .A3(n643), .A4(
        \data_i[12][7] ), .Y(n597) );
  AO22X1_RVT U677 ( .A1(n650), .A2(\data_i[2][7] ), .A3(n649), .A4(
        \data_i[3][7] ), .Y(n604) );
  AO22X1_RVT U678 ( .A1(n652), .A2(\data_i[1][7] ), .A3(n651), .A4(
        \data_i[0][7] ), .Y(n603) );
  AO22X1_RVT U679 ( .A1(n654), .A2(\data_i[6][7] ), .A3(n653), .A4(
        \data_i[7][7] ), .Y(n602) );
  AO22X1_RVT U680 ( .A1(n656), .A2(\data_i[5][7] ), .A3(n655), .A4(
        \data_i[4][7] ), .Y(n601) );
  AO22X1_RVT U681 ( .A1(n662), .A2(\data_i[26][7] ), .A3(n661), .A4(
        \data_i[27][7] ), .Y(n608) );
  AO22X1_RVT U682 ( .A1(n664), .A2(\data_i[25][7] ), .A3(n663), .A4(
        \data_i[24][7] ), .Y(n607) );
  AO22X1_RVT U683 ( .A1(n666), .A2(\data_i[30][7] ), .A3(n665), .A4(
        \data_i[31][7] ), .Y(n606) );
  AO22X1_RVT U684 ( .A1(n668), .A2(\data_i[29][7] ), .A3(n667), .A4(
        \data_i[28][7] ), .Y(n605) );
  AO22X1_RVT U685 ( .A1(n674), .A2(\data_i[18][7] ), .A3(n673), .A4(
        \data_i[19][7] ), .Y(n612) );
  AO22X1_RVT U686 ( .A1(n676), .A2(\data_i[17][7] ), .A3(n675), .A4(
        \data_i[16][7] ), .Y(n611) );
  AO22X1_RVT U687 ( .A1(n678), .A2(\data_i[22][7] ), .A3(n677), .A4(
        \data_i[23][7] ), .Y(n610) );
  AO22X1_RVT U688 ( .A1(n680), .A2(\data_i[21][7] ), .A3(n679), .A4(
        \data_i[20][7] ), .Y(n609) );
  AO22X1_RVT U689 ( .A1(n638), .A2(\data_i[10][8] ), .A3(n637), .A4(
        \data_i[11][8] ), .Y(n620) );
  AO22X1_RVT U690 ( .A1(n640), .A2(\data_i[9][8] ), .A3(n639), .A4(
        \data_i[8][8] ), .Y(n619) );
  AO22X1_RVT U691 ( .A1(n642), .A2(\data_i[14][8] ), .A3(n641), .A4(
        \data_i[15][8] ), .Y(n618) );
  AO22X1_RVT U692 ( .A1(n644), .A2(\data_i[13][8] ), .A3(n643), .A4(
        \data_i[12][8] ), .Y(n617) );
  AO22X1_RVT U693 ( .A1(n650), .A2(\data_i[2][8] ), .A3(n649), .A4(
        \data_i[3][8] ), .Y(n624) );
  AO22X1_RVT U694 ( .A1(n652), .A2(\data_i[1][8] ), .A3(n651), .A4(
        \data_i[0][8] ), .Y(n623) );
  AO22X1_RVT U695 ( .A1(n654), .A2(\data_i[6][8] ), .A3(n653), .A4(
        \data_i[7][8] ), .Y(n622) );
  AO22X1_RVT U696 ( .A1(n656), .A2(\data_i[5][8] ), .A3(n655), .A4(
        \data_i[4][8] ), .Y(n621) );
  AO22X1_RVT U697 ( .A1(n662), .A2(\data_i[26][8] ), .A3(n661), .A4(
        \data_i[27][8] ), .Y(n628) );
  AO22X1_RVT U698 ( .A1(n664), .A2(\data_i[25][8] ), .A3(n663), .A4(
        \data_i[24][8] ), .Y(n627) );
  AO22X1_RVT U699 ( .A1(n666), .A2(\data_i[30][8] ), .A3(n665), .A4(
        \data_i[31][8] ), .Y(n626) );
  AO22X1_RVT U700 ( .A1(n668), .A2(\data_i[29][8] ), .A3(n667), .A4(
        \data_i[28][8] ), .Y(n625) );
  AO22X1_RVT U701 ( .A1(n674), .A2(\data_i[18][8] ), .A3(n673), .A4(
        \data_i[19][8] ), .Y(n632) );
  AO22X1_RVT U702 ( .A1(n676), .A2(\data_i[17][8] ), .A3(n675), .A4(
        \data_i[16][8] ), .Y(n631) );
  AO22X1_RVT U703 ( .A1(n678), .A2(\data_i[22][8] ), .A3(n677), .A4(
        \data_i[23][8] ), .Y(n630) );
  AO22X1_RVT U704 ( .A1(n680), .A2(\data_i[21][8] ), .A3(n679), .A4(
        \data_i[20][8] ), .Y(n629) );
  AO22X1_RVT U705 ( .A1(n638), .A2(\data_i[10][9] ), .A3(n637), .A4(
        \data_i[11][9] ), .Y(n648) );
  AO22X1_RVT U706 ( .A1(n640), .A2(\data_i[9][9] ), .A3(n639), .A4(
        \data_i[8][9] ), .Y(n647) );
  AO22X1_RVT U707 ( .A1(n642), .A2(\data_i[14][9] ), .A3(n641), .A4(
        \data_i[15][9] ), .Y(n646) );
  AO22X1_RVT U708 ( .A1(n644), .A2(\data_i[13][9] ), .A3(n643), .A4(
        \data_i[12][9] ), .Y(n645) );
  AO22X1_RVT U709 ( .A1(n650), .A2(\data_i[2][9] ), .A3(n649), .A4(
        \data_i[3][9] ), .Y(n660) );
  AO22X1_RVT U710 ( .A1(n652), .A2(\data_i[1][9] ), .A3(n651), .A4(
        \data_i[0][9] ), .Y(n659) );
  AO22X1_RVT U711 ( .A1(n654), .A2(\data_i[6][9] ), .A3(n653), .A4(
        \data_i[7][9] ), .Y(n658) );
  AO22X1_RVT U712 ( .A1(n656), .A2(\data_i[5][9] ), .A3(n655), .A4(
        \data_i[4][9] ), .Y(n657) );
  AO22X1_RVT U713 ( .A1(n662), .A2(\data_i[26][9] ), .A3(n661), .A4(
        \data_i[27][9] ), .Y(n672) );
  AO22X1_RVT U714 ( .A1(n664), .A2(\data_i[25][9] ), .A3(n663), .A4(
        \data_i[24][9] ), .Y(n671) );
  AO22X1_RVT U715 ( .A1(n666), .A2(\data_i[30][9] ), .A3(n665), .A4(
        \data_i[31][9] ), .Y(n670) );
  AO22X1_RVT U716 ( .A1(n668), .A2(\data_i[29][9] ), .A3(n667), .A4(
        \data_i[28][9] ), .Y(n669) );
  AO22X1_RVT U717 ( .A1(n674), .A2(\data_i[18][9] ), .A3(n673), .A4(
        \data_i[19][9] ), .Y(n684) );
  AO22X1_RVT U718 ( .A1(n676), .A2(\data_i[17][9] ), .A3(n675), .A4(
        \data_i[16][9] ), .Y(n683) );
  AO22X1_RVT U719 ( .A1(n678), .A2(\data_i[22][9] ), .A3(n677), .A4(
        \data_i[23][9] ), .Y(n682) );
  AO22X1_RVT U720 ( .A1(n680), .A2(\data_i[21][9] ), .A3(n679), .A4(
        \data_i[20][9] ), .Y(n681) );
endmodule


module cam ( reset, clk, read, read_index, write, write_index, write_data, 
        search, search_data, read_valid, read_value, search_valid, 
        search_index );
  input [4:0] read_index;
  input [4:0] write_index;
  input [31:0] write_data;
  input [31:0] search_data;
  output [31:0] read_value;
  output [4:0] search_index;
  input reset, clk, read, write, search;
  output read_valid, search_valid;
  wire   \read_value_mux[31][31] , \read_value_mux[31][30] ,
         \read_value_mux[31][29] , \read_value_mux[31][28] ,
         \read_value_mux[31][27] , \read_value_mux[31][26] ,
         \read_value_mux[31][25] , \read_value_mux[31][24] ,
         \read_value_mux[31][23] , \read_value_mux[31][22] ,
         \read_value_mux[31][21] , \read_value_mux[31][20] ,
         \read_value_mux[31][19] , \read_value_mux[31][18] ,
         \read_value_mux[31][17] , \read_value_mux[31][16] ,
         \read_value_mux[31][15] , \read_value_mux[31][14] ,
         \read_value_mux[31][13] , \read_value_mux[31][12] ,
         \read_value_mux[31][11] , \read_value_mux[31][10] ,
         \read_value_mux[31][9] , \read_value_mux[31][8] ,
         \read_value_mux[31][7] , \read_value_mux[31][6] ,
         \read_value_mux[31][5] , \read_value_mux[31][4] ,
         \read_value_mux[31][3] , \read_value_mux[31][2] ,
         \read_value_mux[31][1] , \read_value_mux[31][0] ,
         \read_value_mux[30][31] , \read_value_mux[30][30] ,
         \read_value_mux[30][29] , \read_value_mux[30][28] ,
         \read_value_mux[30][27] , \read_value_mux[30][26] ,
         \read_value_mux[30][25] , \read_value_mux[30][24] ,
         \read_value_mux[30][23] , \read_value_mux[30][22] ,
         \read_value_mux[30][21] , \read_value_mux[30][20] ,
         \read_value_mux[30][19] , \read_value_mux[30][18] ,
         \read_value_mux[30][17] , \read_value_mux[30][16] ,
         \read_value_mux[30][15] , \read_value_mux[30][14] ,
         \read_value_mux[30][13] , \read_value_mux[30][12] ,
         \read_value_mux[30][11] , \read_value_mux[30][10] ,
         \read_value_mux[30][9] , \read_value_mux[30][8] ,
         \read_value_mux[30][7] , \read_value_mux[30][6] ,
         \read_value_mux[30][5] , \read_value_mux[30][4] ,
         \read_value_mux[30][3] , \read_value_mux[30][2] ,
         \read_value_mux[30][1] , \read_value_mux[30][0] ,
         \read_value_mux[29][31] , \read_value_mux[29][30] ,
         \read_value_mux[29][29] , \read_value_mux[29][28] ,
         \read_value_mux[29][27] , \read_value_mux[29][26] ,
         \read_value_mux[29][25] , \read_value_mux[29][24] ,
         \read_value_mux[29][23] , \read_value_mux[29][22] ,
         \read_value_mux[29][21] , \read_value_mux[29][20] ,
         \read_value_mux[29][19] , \read_value_mux[29][18] ,
         \read_value_mux[29][17] , \read_value_mux[29][16] ,
         \read_value_mux[29][15] , \read_value_mux[29][14] ,
         \read_value_mux[29][13] , \read_value_mux[29][12] ,
         \read_value_mux[29][11] , \read_value_mux[29][10] ,
         \read_value_mux[29][9] , \read_value_mux[29][8] ,
         \read_value_mux[29][7] , \read_value_mux[29][6] ,
         \read_value_mux[29][5] , \read_value_mux[29][4] ,
         \read_value_mux[29][3] , \read_value_mux[29][2] ,
         \read_value_mux[29][1] , \read_value_mux[29][0] ,
         \read_value_mux[28][31] , \read_value_mux[28][30] ,
         \read_value_mux[28][29] , \read_value_mux[28][28] ,
         \read_value_mux[28][27] , \read_value_mux[28][26] ,
         \read_value_mux[28][25] , \read_value_mux[28][24] ,
         \read_value_mux[28][23] , \read_value_mux[28][22] ,
         \read_value_mux[28][21] , \read_value_mux[28][20] ,
         \read_value_mux[28][19] , \read_value_mux[28][18] ,
         \read_value_mux[28][17] , \read_value_mux[28][16] ,
         \read_value_mux[28][15] , \read_value_mux[28][14] ,
         \read_value_mux[28][13] , \read_value_mux[28][12] ,
         \read_value_mux[28][11] , \read_value_mux[28][10] ,
         \read_value_mux[28][9] , \read_value_mux[28][8] ,
         \read_value_mux[28][7] , \read_value_mux[28][6] ,
         \read_value_mux[28][5] , \read_value_mux[28][4] ,
         \read_value_mux[28][3] , \read_value_mux[28][2] ,
         \read_value_mux[28][1] , \read_value_mux[28][0] ,
         \read_value_mux[27][31] , \read_value_mux[27][30] ,
         \read_value_mux[27][29] , \read_value_mux[27][28] ,
         \read_value_mux[27][27] , \read_value_mux[27][26] ,
         \read_value_mux[27][25] , \read_value_mux[27][24] ,
         \read_value_mux[27][23] , \read_value_mux[27][22] ,
         \read_value_mux[27][21] , \read_value_mux[27][20] ,
         \read_value_mux[27][19] , \read_value_mux[27][18] ,
         \read_value_mux[27][17] , \read_value_mux[27][16] ,
         \read_value_mux[27][15] , \read_value_mux[27][14] ,
         \read_value_mux[27][13] , \read_value_mux[27][12] ,
         \read_value_mux[27][11] , \read_value_mux[27][10] ,
         \read_value_mux[27][9] , \read_value_mux[27][8] ,
         \read_value_mux[27][7] , \read_value_mux[27][6] ,
         \read_value_mux[27][5] , \read_value_mux[27][4] ,
         \read_value_mux[27][3] , \read_value_mux[27][2] ,
         \read_value_mux[27][1] , \read_value_mux[27][0] ,
         \read_value_mux[26][31] , \read_value_mux[26][30] ,
         \read_value_mux[26][29] , \read_value_mux[26][28] ,
         \read_value_mux[26][27] , \read_value_mux[26][26] ,
         \read_value_mux[26][25] , \read_value_mux[26][24] ,
         \read_value_mux[26][23] , \read_value_mux[26][22] ,
         \read_value_mux[26][21] , \read_value_mux[26][20] ,
         \read_value_mux[26][19] , \read_value_mux[26][18] ,
         \read_value_mux[26][17] , \read_value_mux[26][16] ,
         \read_value_mux[26][15] , \read_value_mux[26][14] ,
         \read_value_mux[26][13] , \read_value_mux[26][12] ,
         \read_value_mux[26][11] , \read_value_mux[26][10] ,
         \read_value_mux[26][9] , \read_value_mux[26][8] ,
         \read_value_mux[26][7] , \read_value_mux[26][6] ,
         \read_value_mux[26][5] , \read_value_mux[26][4] ,
         \read_value_mux[26][3] , \read_value_mux[26][2] ,
         \read_value_mux[26][1] , \read_value_mux[26][0] ,
         \read_value_mux[25][31] , \read_value_mux[25][30] ,
         \read_value_mux[25][29] , \read_value_mux[25][28] ,
         \read_value_mux[25][27] , \read_value_mux[25][26] ,
         \read_value_mux[25][25] , \read_value_mux[25][24] ,
         \read_value_mux[25][23] , \read_value_mux[25][22] ,
         \read_value_mux[25][21] , \read_value_mux[25][20] ,
         \read_value_mux[25][19] , \read_value_mux[25][18] ,
         \read_value_mux[25][17] , \read_value_mux[25][16] ,
         \read_value_mux[25][15] , \read_value_mux[25][14] ,
         \read_value_mux[25][13] , \read_value_mux[25][12] ,
         \read_value_mux[25][11] , \read_value_mux[25][10] ,
         \read_value_mux[25][9] , \read_value_mux[25][8] ,
         \read_value_mux[25][7] , \read_value_mux[25][6] ,
         \read_value_mux[25][5] , \read_value_mux[25][4] ,
         \read_value_mux[25][3] , \read_value_mux[25][2] ,
         \read_value_mux[25][1] , \read_value_mux[25][0] ,
         \read_value_mux[24][31] , \read_value_mux[24][30] ,
         \read_value_mux[24][29] , \read_value_mux[24][28] ,
         \read_value_mux[24][27] , \read_value_mux[24][26] ,
         \read_value_mux[24][25] , \read_value_mux[24][24] ,
         \read_value_mux[24][23] , \read_value_mux[24][22] ,
         \read_value_mux[24][21] , \read_value_mux[24][20] ,
         \read_value_mux[24][19] , \read_value_mux[24][18] ,
         \read_value_mux[24][17] , \read_value_mux[24][16] ,
         \read_value_mux[24][15] , \read_value_mux[24][14] ,
         \read_value_mux[24][13] , \read_value_mux[24][12] ,
         \read_value_mux[24][11] , \read_value_mux[24][10] ,
         \read_value_mux[24][9] , \read_value_mux[24][8] ,
         \read_value_mux[24][7] , \read_value_mux[24][6] ,
         \read_value_mux[24][5] , \read_value_mux[24][4] ,
         \read_value_mux[24][3] , \read_value_mux[24][2] ,
         \read_value_mux[24][1] , \read_value_mux[24][0] ,
         \read_value_mux[23][31] , \read_value_mux[23][30] ,
         \read_value_mux[23][29] , \read_value_mux[23][28] ,
         \read_value_mux[23][27] , \read_value_mux[23][26] ,
         \read_value_mux[23][25] , \read_value_mux[23][24] ,
         \read_value_mux[23][23] , \read_value_mux[23][22] ,
         \read_value_mux[23][21] , \read_value_mux[23][20] ,
         \read_value_mux[23][19] , \read_value_mux[23][18] ,
         \read_value_mux[23][17] , \read_value_mux[23][16] ,
         \read_value_mux[23][15] , \read_value_mux[23][14] ,
         \read_value_mux[23][13] , \read_value_mux[23][12] ,
         \read_value_mux[23][11] , \read_value_mux[23][10] ,
         \read_value_mux[23][9] , \read_value_mux[23][8] ,
         \read_value_mux[23][7] , \read_value_mux[23][6] ,
         \read_value_mux[23][5] , \read_value_mux[23][4] ,
         \read_value_mux[23][3] , \read_value_mux[23][2] ,
         \read_value_mux[23][1] , \read_value_mux[23][0] ,
         \read_value_mux[22][31] , \read_value_mux[22][30] ,
         \read_value_mux[22][29] , \read_value_mux[22][28] ,
         \read_value_mux[22][27] , \read_value_mux[22][26] ,
         \read_value_mux[22][25] , \read_value_mux[22][24] ,
         \read_value_mux[22][23] , \read_value_mux[22][22] ,
         \read_value_mux[22][21] , \read_value_mux[22][20] ,
         \read_value_mux[22][19] , \read_value_mux[22][18] ,
         \read_value_mux[22][17] , \read_value_mux[22][16] ,
         \read_value_mux[22][15] , \read_value_mux[22][14] ,
         \read_value_mux[22][13] , \read_value_mux[22][12] ,
         \read_value_mux[22][11] , \read_value_mux[22][10] ,
         \read_value_mux[22][9] , \read_value_mux[22][8] ,
         \read_value_mux[22][7] , \read_value_mux[22][6] ,
         \read_value_mux[22][5] , \read_value_mux[22][4] ,
         \read_value_mux[22][3] , \read_value_mux[22][2] ,
         \read_value_mux[22][1] , \read_value_mux[22][0] ,
         \read_value_mux[21][31] , \read_value_mux[21][30] ,
         \read_value_mux[21][29] , \read_value_mux[21][28] ,
         \read_value_mux[21][27] , \read_value_mux[21][26] ,
         \read_value_mux[21][25] , \read_value_mux[21][24] ,
         \read_value_mux[21][23] , \read_value_mux[21][22] ,
         \read_value_mux[21][21] , \read_value_mux[21][20] ,
         \read_value_mux[21][19] , \read_value_mux[21][18] ,
         \read_value_mux[21][17] , \read_value_mux[21][16] ,
         \read_value_mux[21][15] , \read_value_mux[21][14] ,
         \read_value_mux[21][13] , \read_value_mux[21][12] ,
         \read_value_mux[21][11] , \read_value_mux[21][10] ,
         \read_value_mux[21][9] , \read_value_mux[21][8] ,
         \read_value_mux[21][7] , \read_value_mux[21][6] ,
         \read_value_mux[21][5] , \read_value_mux[21][4] ,
         \read_value_mux[21][3] , \read_value_mux[21][2] ,
         \read_value_mux[21][1] , \read_value_mux[21][0] ,
         \read_value_mux[20][31] , \read_value_mux[20][30] ,
         \read_value_mux[20][29] , \read_value_mux[20][28] ,
         \read_value_mux[20][27] , \read_value_mux[20][26] ,
         \read_value_mux[20][25] , \read_value_mux[20][24] ,
         \read_value_mux[20][23] , \read_value_mux[20][22] ,
         \read_value_mux[20][21] , \read_value_mux[20][20] ,
         \read_value_mux[20][19] , \read_value_mux[20][18] ,
         \read_value_mux[20][17] , \read_value_mux[20][16] ,
         \read_value_mux[20][15] , \read_value_mux[20][14] ,
         \read_value_mux[20][13] , \read_value_mux[20][12] ,
         \read_value_mux[20][11] , \read_value_mux[20][10] ,
         \read_value_mux[20][9] , \read_value_mux[20][8] ,
         \read_value_mux[20][7] , \read_value_mux[20][6] ,
         \read_value_mux[20][5] , \read_value_mux[20][4] ,
         \read_value_mux[20][3] , \read_value_mux[20][2] ,
         \read_value_mux[20][1] , \read_value_mux[20][0] ,
         \read_value_mux[19][31] , \read_value_mux[19][30] ,
         \read_value_mux[19][29] , \read_value_mux[19][28] ,
         \read_value_mux[19][27] , \read_value_mux[19][26] ,
         \read_value_mux[19][25] , \read_value_mux[19][24] ,
         \read_value_mux[19][23] , \read_value_mux[19][22] ,
         \read_value_mux[19][21] , \read_value_mux[19][20] ,
         \read_value_mux[19][19] , \read_value_mux[19][18] ,
         \read_value_mux[19][17] , \read_value_mux[19][16] ,
         \read_value_mux[19][15] , \read_value_mux[19][14] ,
         \read_value_mux[19][13] , \read_value_mux[19][12] ,
         \read_value_mux[19][11] , \read_value_mux[19][10] ,
         \read_value_mux[19][9] , \read_value_mux[19][8] ,
         \read_value_mux[19][7] , \read_value_mux[19][6] ,
         \read_value_mux[19][5] , \read_value_mux[19][4] ,
         \read_value_mux[19][3] , \read_value_mux[19][2] ,
         \read_value_mux[19][1] , \read_value_mux[19][0] ,
         \read_value_mux[18][31] , \read_value_mux[18][30] ,
         \read_value_mux[18][29] , \read_value_mux[18][28] ,
         \read_value_mux[18][27] , \read_value_mux[18][26] ,
         \read_value_mux[18][25] , \read_value_mux[18][24] ,
         \read_value_mux[18][23] , \read_value_mux[18][22] ,
         \read_value_mux[18][21] , \read_value_mux[18][20] ,
         \read_value_mux[18][19] , \read_value_mux[18][18] ,
         \read_value_mux[18][17] , \read_value_mux[18][16] ,
         \read_value_mux[18][15] , \read_value_mux[18][14] ,
         \read_value_mux[18][13] , \read_value_mux[18][12] ,
         \read_value_mux[18][11] , \read_value_mux[18][10] ,
         \read_value_mux[18][9] , \read_value_mux[18][8] ,
         \read_value_mux[18][7] , \read_value_mux[18][6] ,
         \read_value_mux[18][5] , \read_value_mux[18][4] ,
         \read_value_mux[18][3] , \read_value_mux[18][2] ,
         \read_value_mux[18][1] , \read_value_mux[18][0] ,
         \read_value_mux[17][31] , \read_value_mux[17][30] ,
         \read_value_mux[17][29] , \read_value_mux[17][28] ,
         \read_value_mux[17][27] , \read_value_mux[17][26] ,
         \read_value_mux[17][25] , \read_value_mux[17][24] ,
         \read_value_mux[17][23] , \read_value_mux[17][22] ,
         \read_value_mux[17][21] , \read_value_mux[17][20] ,
         \read_value_mux[17][19] , \read_value_mux[17][18] ,
         \read_value_mux[17][17] , \read_value_mux[17][16] ,
         \read_value_mux[17][15] , \read_value_mux[17][14] ,
         \read_value_mux[17][13] , \read_value_mux[17][12] ,
         \read_value_mux[17][11] , \read_value_mux[17][10] ,
         \read_value_mux[17][9] , \read_value_mux[17][8] ,
         \read_value_mux[17][7] , \read_value_mux[17][6] ,
         \read_value_mux[17][5] , \read_value_mux[17][4] ,
         \read_value_mux[17][3] , \read_value_mux[17][2] ,
         \read_value_mux[17][1] , \read_value_mux[17][0] ,
         \read_value_mux[16][31] , \read_value_mux[16][30] ,
         \read_value_mux[16][29] , \read_value_mux[16][28] ,
         \read_value_mux[16][27] , \read_value_mux[16][26] ,
         \read_value_mux[16][25] , \read_value_mux[16][24] ,
         \read_value_mux[16][23] , \read_value_mux[16][22] ,
         \read_value_mux[16][21] , \read_value_mux[16][20] ,
         \read_value_mux[16][19] , \read_value_mux[16][18] ,
         \read_value_mux[16][17] , \read_value_mux[16][16] ,
         \read_value_mux[16][15] , \read_value_mux[16][14] ,
         \read_value_mux[16][13] , \read_value_mux[16][12] ,
         \read_value_mux[16][11] , \read_value_mux[16][10] ,
         \read_value_mux[16][9] , \read_value_mux[16][8] ,
         \read_value_mux[16][7] , \read_value_mux[16][6] ,
         \read_value_mux[16][5] , \read_value_mux[16][4] ,
         \read_value_mux[16][3] , \read_value_mux[16][2] ,
         \read_value_mux[16][1] , \read_value_mux[16][0] ,
         \read_value_mux[15][31] , \read_value_mux[15][30] ,
         \read_value_mux[15][29] , \read_value_mux[15][28] ,
         \read_value_mux[15][27] , \read_value_mux[15][26] ,
         \read_value_mux[15][25] , \read_value_mux[15][24] ,
         \read_value_mux[15][23] , \read_value_mux[15][22] ,
         \read_value_mux[15][21] , \read_value_mux[15][20] ,
         \read_value_mux[15][19] , \read_value_mux[15][18] ,
         \read_value_mux[15][17] , \read_value_mux[15][16] ,
         \read_value_mux[15][15] , \read_value_mux[15][14] ,
         \read_value_mux[15][13] , \read_value_mux[15][12] ,
         \read_value_mux[15][11] , \read_value_mux[15][10] ,
         \read_value_mux[15][9] , \read_value_mux[15][8] ,
         \read_value_mux[15][7] , \read_value_mux[15][6] ,
         \read_value_mux[15][5] , \read_value_mux[15][4] ,
         \read_value_mux[15][3] , \read_value_mux[15][2] ,
         \read_value_mux[15][1] , \read_value_mux[15][0] ,
         \read_value_mux[14][31] , \read_value_mux[14][30] ,
         \read_value_mux[14][29] , \read_value_mux[14][28] ,
         \read_value_mux[14][27] , \read_value_mux[14][26] ,
         \read_value_mux[14][25] , \read_value_mux[14][24] ,
         \read_value_mux[14][23] , \read_value_mux[14][22] ,
         \read_value_mux[14][21] , \read_value_mux[14][20] ,
         \read_value_mux[14][19] , \read_value_mux[14][18] ,
         \read_value_mux[14][17] , \read_value_mux[14][16] ,
         \read_value_mux[14][15] , \read_value_mux[14][14] ,
         \read_value_mux[14][13] , \read_value_mux[14][12] ,
         \read_value_mux[14][11] , \read_value_mux[14][10] ,
         \read_value_mux[14][9] , \read_value_mux[14][8] ,
         \read_value_mux[14][7] , \read_value_mux[14][6] ,
         \read_value_mux[14][5] , \read_value_mux[14][4] ,
         \read_value_mux[14][3] , \read_value_mux[14][2] ,
         \read_value_mux[14][1] , \read_value_mux[14][0] ,
         \read_value_mux[13][31] , \read_value_mux[13][30] ,
         \read_value_mux[13][29] , \read_value_mux[13][28] ,
         \read_value_mux[13][27] , \read_value_mux[13][26] ,
         \read_value_mux[13][25] , \read_value_mux[13][24] ,
         \read_value_mux[13][23] , \read_value_mux[13][22] ,
         \read_value_mux[13][21] , \read_value_mux[13][20] ,
         \read_value_mux[13][19] , \read_value_mux[13][18] ,
         \read_value_mux[13][17] , \read_value_mux[13][16] ,
         \read_value_mux[13][15] , \read_value_mux[13][14] ,
         \read_value_mux[13][13] , \read_value_mux[13][12] ,
         \read_value_mux[13][11] , \read_value_mux[13][10] ,
         \read_value_mux[13][9] , \read_value_mux[13][8] ,
         \read_value_mux[13][7] , \read_value_mux[13][6] ,
         \read_value_mux[13][5] , \read_value_mux[13][4] ,
         \read_value_mux[13][3] , \read_value_mux[13][2] ,
         \read_value_mux[13][1] , \read_value_mux[13][0] ,
         \read_value_mux[12][31] , \read_value_mux[12][30] ,
         \read_value_mux[12][29] , \read_value_mux[12][28] ,
         \read_value_mux[12][27] , \read_value_mux[12][26] ,
         \read_value_mux[12][25] , \read_value_mux[12][24] ,
         \read_value_mux[12][23] , \read_value_mux[12][22] ,
         \read_value_mux[12][21] , \read_value_mux[12][20] ,
         \read_value_mux[12][19] , \read_value_mux[12][18] ,
         \read_value_mux[12][17] , \read_value_mux[12][16] ,
         \read_value_mux[12][15] , \read_value_mux[12][14] ,
         \read_value_mux[12][13] , \read_value_mux[12][12] ,
         \read_value_mux[12][11] , \read_value_mux[12][10] ,
         \read_value_mux[12][9] , \read_value_mux[12][8] ,
         \read_value_mux[12][7] , \read_value_mux[12][6] ,
         \read_value_mux[12][5] , \read_value_mux[12][4] ,
         \read_value_mux[12][3] , \read_value_mux[12][2] ,
         \read_value_mux[12][1] , \read_value_mux[12][0] ,
         \read_value_mux[11][31] , \read_value_mux[11][30] ,
         \read_value_mux[11][29] , \read_value_mux[11][28] ,
         \read_value_mux[11][27] , \read_value_mux[11][26] ,
         \read_value_mux[11][25] , \read_value_mux[11][24] ,
         \read_value_mux[11][23] , \read_value_mux[11][22] ,
         \read_value_mux[11][21] , \read_value_mux[11][20] ,
         \read_value_mux[11][19] , \read_value_mux[11][18] ,
         \read_value_mux[11][17] , \read_value_mux[11][16] ,
         \read_value_mux[11][15] , \read_value_mux[11][14] ,
         \read_value_mux[11][13] , \read_value_mux[11][12] ,
         \read_value_mux[11][11] , \read_value_mux[11][10] ,
         \read_value_mux[11][9] , \read_value_mux[11][8] ,
         \read_value_mux[11][7] , \read_value_mux[11][6] ,
         \read_value_mux[11][5] , \read_value_mux[11][4] ,
         \read_value_mux[11][3] , \read_value_mux[11][2] ,
         \read_value_mux[11][1] , \read_value_mux[11][0] ,
         \read_value_mux[10][31] , \read_value_mux[10][30] ,
         \read_value_mux[10][29] , \read_value_mux[10][28] ,
         \read_value_mux[10][27] , \read_value_mux[10][26] ,
         \read_value_mux[10][25] , \read_value_mux[10][24] ,
         \read_value_mux[10][23] , \read_value_mux[10][22] ,
         \read_value_mux[10][21] , \read_value_mux[10][20] ,
         \read_value_mux[10][19] , \read_value_mux[10][18] ,
         \read_value_mux[10][17] , \read_value_mux[10][16] ,
         \read_value_mux[10][15] , \read_value_mux[10][14] ,
         \read_value_mux[10][13] , \read_value_mux[10][12] ,
         \read_value_mux[10][11] , \read_value_mux[10][10] ,
         \read_value_mux[10][9] , \read_value_mux[10][8] ,
         \read_value_mux[10][7] , \read_value_mux[10][6] ,
         \read_value_mux[10][5] , \read_value_mux[10][4] ,
         \read_value_mux[10][3] , \read_value_mux[10][2] ,
         \read_value_mux[10][1] , \read_value_mux[10][0] ,
         \read_value_mux[9][31] , \read_value_mux[9][30] ,
         \read_value_mux[9][29] , \read_value_mux[9][28] ,
         \read_value_mux[9][27] , \read_value_mux[9][26] ,
         \read_value_mux[9][25] , \read_value_mux[9][24] ,
         \read_value_mux[9][23] , \read_value_mux[9][22] ,
         \read_value_mux[9][21] , \read_value_mux[9][20] ,
         \read_value_mux[9][19] , \read_value_mux[9][18] ,
         \read_value_mux[9][17] , \read_value_mux[9][16] ,
         \read_value_mux[9][15] , \read_value_mux[9][14] ,
         \read_value_mux[9][13] , \read_value_mux[9][12] ,
         \read_value_mux[9][11] , \read_value_mux[9][10] ,
         \read_value_mux[9][9] , \read_value_mux[9][8] ,
         \read_value_mux[9][7] , \read_value_mux[9][6] ,
         \read_value_mux[9][5] , \read_value_mux[9][4] ,
         \read_value_mux[9][3] , \read_value_mux[9][2] ,
         \read_value_mux[9][1] , \read_value_mux[9][0] ,
         \read_value_mux[8][31] , \read_value_mux[8][30] ,
         \read_value_mux[8][29] , \read_value_mux[8][28] ,
         \read_value_mux[8][27] , \read_value_mux[8][26] ,
         \read_value_mux[8][25] , \read_value_mux[8][24] ,
         \read_value_mux[8][23] , \read_value_mux[8][22] ,
         \read_value_mux[8][21] , \read_value_mux[8][20] ,
         \read_value_mux[8][19] , \read_value_mux[8][18] ,
         \read_value_mux[8][17] , \read_value_mux[8][16] ,
         \read_value_mux[8][15] , \read_value_mux[8][14] ,
         \read_value_mux[8][13] , \read_value_mux[8][12] ,
         \read_value_mux[8][11] , \read_value_mux[8][10] ,
         \read_value_mux[8][9] , \read_value_mux[8][8] ,
         \read_value_mux[8][7] , \read_value_mux[8][6] ,
         \read_value_mux[8][5] , \read_value_mux[8][4] ,
         \read_value_mux[8][3] , \read_value_mux[8][2] ,
         \read_value_mux[8][1] , \read_value_mux[8][0] ,
         \read_value_mux[7][31] , \read_value_mux[7][30] ,
         \read_value_mux[7][29] , \read_value_mux[7][28] ,
         \read_value_mux[7][27] , \read_value_mux[7][26] ,
         \read_value_mux[7][25] , \read_value_mux[7][24] ,
         \read_value_mux[7][23] , \read_value_mux[7][22] ,
         \read_value_mux[7][21] , \read_value_mux[7][20] ,
         \read_value_mux[7][19] , \read_value_mux[7][18] ,
         \read_value_mux[7][17] , \read_value_mux[7][16] ,
         \read_value_mux[7][15] , \read_value_mux[7][14] ,
         \read_value_mux[7][13] , \read_value_mux[7][12] ,
         \read_value_mux[7][11] , \read_value_mux[7][10] ,
         \read_value_mux[7][9] , \read_value_mux[7][8] ,
         \read_value_mux[7][7] , \read_value_mux[7][6] ,
         \read_value_mux[7][5] , \read_value_mux[7][4] ,
         \read_value_mux[7][3] , \read_value_mux[7][2] ,
         \read_value_mux[7][1] , \read_value_mux[7][0] ,
         \read_value_mux[6][31] , \read_value_mux[6][30] ,
         \read_value_mux[6][29] , \read_value_mux[6][28] ,
         \read_value_mux[6][27] , \read_value_mux[6][26] ,
         \read_value_mux[6][25] , \read_value_mux[6][24] ,
         \read_value_mux[6][23] , \read_value_mux[6][22] ,
         \read_value_mux[6][21] , \read_value_mux[6][20] ,
         \read_value_mux[6][19] , \read_value_mux[6][18] ,
         \read_value_mux[6][17] , \read_value_mux[6][16] ,
         \read_value_mux[6][15] , \read_value_mux[6][14] ,
         \read_value_mux[6][13] , \read_value_mux[6][12] ,
         \read_value_mux[6][11] , \read_value_mux[6][10] ,
         \read_value_mux[6][9] , \read_value_mux[6][8] ,
         \read_value_mux[6][7] , \read_value_mux[6][6] ,
         \read_value_mux[6][5] , \read_value_mux[6][4] ,
         \read_value_mux[6][3] , \read_value_mux[6][2] ,
         \read_value_mux[6][1] , \read_value_mux[6][0] ,
         \read_value_mux[5][31] , \read_value_mux[5][30] ,
         \read_value_mux[5][29] , \read_value_mux[5][28] ,
         \read_value_mux[5][27] , \read_value_mux[5][26] ,
         \read_value_mux[5][25] , \read_value_mux[5][24] ,
         \read_value_mux[5][23] , \read_value_mux[5][22] ,
         \read_value_mux[5][21] , \read_value_mux[5][20] ,
         \read_value_mux[5][19] , \read_value_mux[5][18] ,
         \read_value_mux[5][17] , \read_value_mux[5][16] ,
         \read_value_mux[5][15] , \read_value_mux[5][14] ,
         \read_value_mux[5][13] , \read_value_mux[5][12] ,
         \read_value_mux[5][11] , \read_value_mux[5][10] ,
         \read_value_mux[5][9] , \read_value_mux[5][8] ,
         \read_value_mux[5][7] , \read_value_mux[5][6] ,
         \read_value_mux[5][5] , \read_value_mux[5][4] ,
         \read_value_mux[5][3] , \read_value_mux[5][2] ,
         \read_value_mux[5][1] , \read_value_mux[5][0] ,
         \read_value_mux[4][31] , \read_value_mux[4][30] ,
         \read_value_mux[4][29] , \read_value_mux[4][28] ,
         \read_value_mux[4][27] , \read_value_mux[4][26] ,
         \read_value_mux[4][25] , \read_value_mux[4][24] ,
         \read_value_mux[4][23] , \read_value_mux[4][22] ,
         \read_value_mux[4][21] , \read_value_mux[4][20] ,
         \read_value_mux[4][19] , \read_value_mux[4][18] ,
         \read_value_mux[4][17] , \read_value_mux[4][16] ,
         \read_value_mux[4][15] , \read_value_mux[4][14] ,
         \read_value_mux[4][13] , \read_value_mux[4][12] ,
         \read_value_mux[4][11] , \read_value_mux[4][10] ,
         \read_value_mux[4][9] , \read_value_mux[4][8] ,
         \read_value_mux[4][7] , \read_value_mux[4][6] ,
         \read_value_mux[4][5] , \read_value_mux[4][4] ,
         \read_value_mux[4][3] , \read_value_mux[4][2] ,
         \read_value_mux[4][1] , \read_value_mux[4][0] ,
         \read_value_mux[3][31] , \read_value_mux[3][30] ,
         \read_value_mux[3][29] , \read_value_mux[3][28] ,
         \read_value_mux[3][27] , \read_value_mux[3][26] ,
         \read_value_mux[3][25] , \read_value_mux[3][24] ,
         \read_value_mux[3][23] , \read_value_mux[3][22] ,
         \read_value_mux[3][21] , \read_value_mux[3][20] ,
         \read_value_mux[3][19] , \read_value_mux[3][18] ,
         \read_value_mux[3][17] , \read_value_mux[3][16] ,
         \read_value_mux[3][15] , \read_value_mux[3][14] ,
         \read_value_mux[3][13] , \read_value_mux[3][12] ,
         \read_value_mux[3][11] , \read_value_mux[3][10] ,
         \read_value_mux[3][9] , \read_value_mux[3][8] ,
         \read_value_mux[3][7] , \read_value_mux[3][6] ,
         \read_value_mux[3][5] , \read_value_mux[3][4] ,
         \read_value_mux[3][3] , \read_value_mux[3][2] ,
         \read_value_mux[3][1] , \read_value_mux[3][0] ,
         \read_value_mux[2][31] , \read_value_mux[2][30] ,
         \read_value_mux[2][29] , \read_value_mux[2][28] ,
         \read_value_mux[2][27] , \read_value_mux[2][26] ,
         \read_value_mux[2][25] , \read_value_mux[2][24] ,
         \read_value_mux[2][23] , \read_value_mux[2][22] ,
         \read_value_mux[2][21] , \read_value_mux[2][20] ,
         \read_value_mux[2][19] , \read_value_mux[2][18] ,
         \read_value_mux[2][17] , \read_value_mux[2][16] ,
         \read_value_mux[2][15] , \read_value_mux[2][14] ,
         \read_value_mux[2][13] , \read_value_mux[2][12] ,
         \read_value_mux[2][11] , \read_value_mux[2][10] ,
         \read_value_mux[2][9] , \read_value_mux[2][8] ,
         \read_value_mux[2][7] , \read_value_mux[2][6] ,
         \read_value_mux[2][5] , \read_value_mux[2][4] ,
         \read_value_mux[2][3] , \read_value_mux[2][2] ,
         \read_value_mux[2][1] , \read_value_mux[2][0] ,
         \read_value_mux[1][31] , \read_value_mux[1][30] ,
         \read_value_mux[1][29] , \read_value_mux[1][28] ,
         \read_value_mux[1][27] , \read_value_mux[1][26] ,
         \read_value_mux[1][25] , \read_value_mux[1][24] ,
         \read_value_mux[1][23] , \read_value_mux[1][22] ,
         \read_value_mux[1][21] , \read_value_mux[1][20] ,
         \read_value_mux[1][19] , \read_value_mux[1][18] ,
         \read_value_mux[1][17] , \read_value_mux[1][16] ,
         \read_value_mux[1][15] , \read_value_mux[1][14] ,
         \read_value_mux[1][13] , \read_value_mux[1][12] ,
         \read_value_mux[1][11] , \read_value_mux[1][10] ,
         \read_value_mux[1][9] , \read_value_mux[1][8] ,
         \read_value_mux[1][7] , \read_value_mux[1][6] ,
         \read_value_mux[1][5] , \read_value_mux[1][4] ,
         \read_value_mux[1][3] , \read_value_mux[1][2] ,
         \read_value_mux[1][1] , \read_value_mux[1][0] ,
         \read_value_mux[0][31] , \read_value_mux[0][30] ,
         \read_value_mux[0][29] , \read_value_mux[0][28] ,
         \read_value_mux[0][27] , \read_value_mux[0][26] ,
         \read_value_mux[0][25] , \read_value_mux[0][24] ,
         \read_value_mux[0][23] , \read_value_mux[0][22] ,
         \read_value_mux[0][21] , \read_value_mux[0][20] ,
         \read_value_mux[0][19] , \read_value_mux[0][18] ,
         \read_value_mux[0][17] , \read_value_mux[0][16] ,
         \read_value_mux[0][15] , \read_value_mux[0][14] ,
         \read_value_mux[0][13] , \read_value_mux[0][12] ,
         \read_value_mux[0][11] , \read_value_mux[0][10] ,
         \read_value_mux[0][9] , \read_value_mux[0][8] ,
         \read_value_mux[0][7] , \read_value_mux[0][6] ,
         \read_value_mux[0][5] , \read_value_mux[0][4] ,
         \read_value_mux[0][3] , \read_value_mux[0][2] ,
         \read_value_mux[0][1] , \read_value_mux[0][0] , \words[31]/valid_o ,
         \words[31]/valid_i , \words[31]/data_i[31] , \words[31]/data_i[30] ,
         \words[31]/data_i[29] , \words[31]/data_i[28] ,
         \words[31]/data_i[27] , \words[31]/data_i[26] ,
         \words[31]/data_i[25] , \words[31]/data_i[24] ,
         \words[31]/data_i[23] , \words[31]/data_i[22] ,
         \words[31]/data_i[21] , \words[31]/data_i[20] ,
         \words[31]/data_i[19] , \words[31]/data_i[18] ,
         \words[31]/data_i[17] , \words[31]/data_i[16] ,
         \words[31]/data_i[15] , \words[31]/data_i[14] ,
         \words[31]/data_i[13] , \words[31]/data_i[12] ,
         \words[31]/data_i[11] , \words[31]/data_i[10] , \words[31]/data_i[9] ,
         \words[31]/data_i[8] , \words[31]/data_i[7] , \words[31]/data_i[6] ,
         \words[31]/data_i[5] , \words[31]/data_i[4] , \words[31]/data_i[3] ,
         \words[31]/data_i[2] , \words[31]/data_i[1] , \words[31]/data_i[0] ,
         \words[0]/valid_o , \words[0]/valid_i , \words[0]/data_i[31] ,
         \words[0]/data_i[30] , \words[0]/data_i[29] , \words[0]/data_i[28] ,
         \words[0]/data_i[27] , \words[0]/data_i[26] , \words[0]/data_i[25] ,
         \words[0]/data_i[24] , \words[0]/data_i[23] , \words[0]/data_i[22] ,
         \words[0]/data_i[21] , \words[0]/data_i[20] , \words[0]/data_i[19] ,
         \words[0]/data_i[18] , \words[0]/data_i[17] , \words[0]/data_i[16] ,
         \words[0]/data_i[15] , \words[0]/data_i[14] , \words[0]/data_i[13] ,
         \words[0]/data_i[12] , \words[0]/data_i[11] , \words[0]/data_i[10] ,
         \words[0]/data_i[9] , \words[0]/data_i[8] , \words[0]/data_i[7] ,
         \words[0]/data_i[6] , \words[0]/data_i[5] , \words[0]/data_i[4] ,
         \words[0]/data_i[3] , \words[0]/data_i[2] , \words[0]/data_i[1] ,
         \words[0]/data_i[0] , \words[1]/valid_o , \words[1]/valid_i ,
         \words[1]/data_i[31] , \words[1]/data_i[30] , \words[1]/data_i[29] ,
         \words[1]/data_i[28] , \words[1]/data_i[27] , \words[1]/data_i[26] ,
         \words[1]/data_i[25] , \words[1]/data_i[24] , \words[1]/data_i[23] ,
         \words[1]/data_i[22] , \words[1]/data_i[21] , \words[1]/data_i[20] ,
         \words[1]/data_i[19] , \words[1]/data_i[18] , \words[1]/data_i[17] ,
         \words[1]/data_i[16] , \words[1]/data_i[15] , \words[1]/data_i[14] ,
         \words[1]/data_i[13] , \words[1]/data_i[12] , \words[1]/data_i[11] ,
         \words[1]/data_i[10] , \words[1]/data_i[9] , \words[1]/data_i[8] ,
         \words[1]/data_i[7] , \words[1]/data_i[6] , \words[1]/data_i[5] ,
         \words[1]/data_i[4] , \words[1]/data_i[3] , \words[1]/data_i[2] ,
         \words[1]/data_i[1] , \words[1]/data_i[0] , \words[2]/valid_o ,
         \words[2]/valid_i , \words[2]/data_i[31] , \words[2]/data_i[30] ,
         \words[2]/data_i[29] , \words[2]/data_i[28] , \words[2]/data_i[27] ,
         \words[2]/data_i[26] , \words[2]/data_i[25] , \words[2]/data_i[24] ,
         \words[2]/data_i[23] , \words[2]/data_i[22] , \words[2]/data_i[21] ,
         \words[2]/data_i[20] , \words[2]/data_i[19] , \words[2]/data_i[18] ,
         \words[2]/data_i[17] , \words[2]/data_i[16] , \words[2]/data_i[15] ,
         \words[2]/data_i[14] , \words[2]/data_i[13] , \words[2]/data_i[12] ,
         \words[2]/data_i[11] , \words[2]/data_i[10] , \words[2]/data_i[9] ,
         \words[2]/data_i[8] , \words[2]/data_i[7] , \words[2]/data_i[6] ,
         \words[2]/data_i[5] , \words[2]/data_i[4] , \words[2]/data_i[3] ,
         \words[2]/data_i[2] , \words[2]/data_i[1] , \words[2]/data_i[0] ,
         \words[3]/valid_o , \words[3]/valid_i , \words[3]/data_i[31] ,
         \words[3]/data_i[30] , \words[3]/data_i[29] , \words[3]/data_i[28] ,
         \words[3]/data_i[27] , \words[3]/data_i[26] , \words[3]/data_i[25] ,
         \words[3]/data_i[24] , \words[3]/data_i[23] , \words[3]/data_i[22] ,
         \words[3]/data_i[21] , \words[3]/data_i[20] , \words[3]/data_i[19] ,
         \words[3]/data_i[18] , \words[3]/data_i[17] , \words[3]/data_i[16] ,
         \words[3]/data_i[15] , \words[3]/data_i[14] , \words[3]/data_i[13] ,
         \words[3]/data_i[12] , \words[3]/data_i[11] , \words[3]/data_i[10] ,
         \words[3]/data_i[9] , \words[3]/data_i[8] , \words[3]/data_i[7] ,
         \words[3]/data_i[6] , \words[3]/data_i[5] , \words[3]/data_i[4] ,
         \words[3]/data_i[3] , \words[3]/data_i[2] , \words[3]/data_i[1] ,
         \words[3]/data_i[0] , \words[4]/valid_o , \words[4]/valid_i ,
         \words[4]/data_i[31] , \words[4]/data_i[30] , \words[4]/data_i[29] ,
         \words[4]/data_i[28] , \words[4]/data_i[27] , \words[4]/data_i[26] ,
         \words[4]/data_i[25] , \words[4]/data_i[24] , \words[4]/data_i[23] ,
         \words[4]/data_i[22] , \words[4]/data_i[21] , \words[4]/data_i[20] ,
         \words[4]/data_i[19] , \words[4]/data_i[18] , \words[4]/data_i[17] ,
         \words[4]/data_i[16] , \words[4]/data_i[15] , \words[4]/data_i[14] ,
         \words[4]/data_i[13] , \words[4]/data_i[12] , \words[4]/data_i[11] ,
         \words[4]/data_i[10] , \words[4]/data_i[9] , \words[4]/data_i[8] ,
         \words[4]/data_i[7] , \words[4]/data_i[6] , \words[4]/data_i[5] ,
         \words[4]/data_i[4] , \words[4]/data_i[3] , \words[4]/data_i[2] ,
         \words[4]/data_i[1] , \words[4]/data_i[0] , \words[5]/valid_o ,
         \words[5]/valid_i , \words[5]/data_i[31] , \words[5]/data_i[30] ,
         \words[5]/data_i[29] , \words[5]/data_i[28] , \words[5]/data_i[27] ,
         \words[5]/data_i[26] , \words[5]/data_i[25] , \words[5]/data_i[24] ,
         \words[5]/data_i[23] , \words[5]/data_i[22] , \words[5]/data_i[21] ,
         \words[5]/data_i[20] , \words[5]/data_i[19] , \words[5]/data_i[18] ,
         \words[5]/data_i[17] , \words[5]/data_i[16] , \words[5]/data_i[15] ,
         \words[5]/data_i[14] , \words[5]/data_i[13] , \words[5]/data_i[12] ,
         \words[5]/data_i[11] , \words[5]/data_i[10] , \words[5]/data_i[9] ,
         \words[5]/data_i[8] , \words[5]/data_i[7] , \words[5]/data_i[6] ,
         \words[5]/data_i[5] , \words[5]/data_i[4] , \words[5]/data_i[3] ,
         \words[5]/data_i[2] , \words[5]/data_i[1] , \words[5]/data_i[0] ,
         \words[6]/valid_o , \words[6]/valid_i , \words[6]/data_i[31] ,
         \words[6]/data_i[30] , \words[6]/data_i[29] , \words[6]/data_i[28] ,
         \words[6]/data_i[27] , \words[6]/data_i[26] , \words[6]/data_i[25] ,
         \words[6]/data_i[24] , \words[6]/data_i[23] , \words[6]/data_i[22] ,
         \words[6]/data_i[21] , \words[6]/data_i[20] , \words[6]/data_i[19] ,
         \words[6]/data_i[18] , \words[6]/data_i[17] , \words[6]/data_i[16] ,
         \words[6]/data_i[15] , \words[6]/data_i[14] , \words[6]/data_i[13] ,
         \words[6]/data_i[12] , \words[6]/data_i[11] , \words[6]/data_i[10] ,
         \words[6]/data_i[9] , \words[6]/data_i[8] , \words[6]/data_i[7] ,
         \words[6]/data_i[6] , \words[6]/data_i[5] , \words[6]/data_i[4] ,
         \words[6]/data_i[3] , \words[6]/data_i[2] , \words[6]/data_i[1] ,
         \words[6]/data_i[0] , \words[7]/valid_o , \words[7]/valid_i ,
         \words[7]/data_i[31] , \words[7]/data_i[30] , \words[7]/data_i[29] ,
         \words[7]/data_i[28] , \words[7]/data_i[27] , \words[7]/data_i[26] ,
         \words[7]/data_i[25] , \words[7]/data_i[24] , \words[7]/data_i[23] ,
         \words[7]/data_i[22] , \words[7]/data_i[21] , \words[7]/data_i[20] ,
         \words[7]/data_i[19] , \words[7]/data_i[18] , \words[7]/data_i[17] ,
         \words[7]/data_i[16] , \words[7]/data_i[15] , \words[7]/data_i[14] ,
         \words[7]/data_i[13] , \words[7]/data_i[12] , \words[7]/data_i[11] ,
         \words[7]/data_i[10] , \words[7]/data_i[9] , \words[7]/data_i[8] ,
         \words[7]/data_i[7] , \words[7]/data_i[6] , \words[7]/data_i[5] ,
         \words[7]/data_i[4] , \words[7]/data_i[3] , \words[7]/data_i[2] ,
         \words[7]/data_i[1] , \words[7]/data_i[0] , \words[8]/valid_o ,
         \words[8]/valid_i , \words[8]/data_i[31] , \words[8]/data_i[30] ,
         \words[8]/data_i[29] , \words[8]/data_i[28] , \words[8]/data_i[27] ,
         \words[8]/data_i[26] , \words[8]/data_i[25] , \words[8]/data_i[24] ,
         \words[8]/data_i[23] , \words[8]/data_i[22] , \words[8]/data_i[21] ,
         \words[8]/data_i[20] , \words[8]/data_i[19] , \words[8]/data_i[18] ,
         \words[8]/data_i[17] , \words[8]/data_i[16] , \words[8]/data_i[15] ,
         \words[8]/data_i[14] , \words[8]/data_i[13] , \words[8]/data_i[12] ,
         \words[8]/data_i[11] , \words[8]/data_i[10] , \words[8]/data_i[9] ,
         \words[8]/data_i[8] , \words[8]/data_i[7] , \words[8]/data_i[6] ,
         \words[8]/data_i[5] , \words[8]/data_i[4] , \words[8]/data_i[3] ,
         \words[8]/data_i[2] , \words[8]/data_i[1] , \words[8]/data_i[0] ,
         \words[9]/valid_o , \words[9]/valid_i , \words[9]/data_i[31] ,
         \words[9]/data_i[30] , \words[9]/data_i[29] , \words[9]/data_i[28] ,
         \words[9]/data_i[27] , \words[9]/data_i[26] , \words[9]/data_i[25] ,
         \words[9]/data_i[24] , \words[9]/data_i[23] , \words[9]/data_i[22] ,
         \words[9]/data_i[21] , \words[9]/data_i[20] , \words[9]/data_i[19] ,
         \words[9]/data_i[18] , \words[9]/data_i[17] , \words[9]/data_i[16] ,
         \words[9]/data_i[15] , \words[9]/data_i[14] , \words[9]/data_i[13] ,
         \words[9]/data_i[12] , \words[9]/data_i[11] , \words[9]/data_i[10] ,
         \words[9]/data_i[9] , \words[9]/data_i[8] , \words[9]/data_i[7] ,
         \words[9]/data_i[6] , \words[9]/data_i[5] , \words[9]/data_i[4] ,
         \words[9]/data_i[3] , \words[9]/data_i[2] , \words[9]/data_i[1] ,
         \words[9]/data_i[0] , \words[10]/valid_o , \words[10]/valid_i ,
         \words[10]/data_i[31] , \words[10]/data_i[30] ,
         \words[10]/data_i[29] , \words[10]/data_i[28] ,
         \words[10]/data_i[27] , \words[10]/data_i[26] ,
         \words[10]/data_i[25] , \words[10]/data_i[24] ,
         \words[10]/data_i[23] , \words[10]/data_i[22] ,
         \words[10]/data_i[21] , \words[10]/data_i[20] ,
         \words[10]/data_i[19] , \words[10]/data_i[18] ,
         \words[10]/data_i[17] , \words[10]/data_i[16] ,
         \words[10]/data_i[15] , \words[10]/data_i[14] ,
         \words[10]/data_i[13] , \words[10]/data_i[12] ,
         \words[10]/data_i[11] , \words[10]/data_i[10] , \words[10]/data_i[9] ,
         \words[10]/data_i[8] , \words[10]/data_i[7] , \words[10]/data_i[6] ,
         \words[10]/data_i[5] , \words[10]/data_i[4] , \words[10]/data_i[3] ,
         \words[10]/data_i[2] , \words[10]/data_i[1] , \words[10]/data_i[0] ,
         \words[11]/valid_o , \words[11]/valid_i , \words[11]/data_i[31] ,
         \words[11]/data_i[30] , \words[11]/data_i[29] ,
         \words[11]/data_i[28] , \words[11]/data_i[27] ,
         \words[11]/data_i[26] , \words[11]/data_i[25] ,
         \words[11]/data_i[24] , \words[11]/data_i[23] ,
         \words[11]/data_i[22] , \words[11]/data_i[21] ,
         \words[11]/data_i[20] , \words[11]/data_i[19] ,
         \words[11]/data_i[18] , \words[11]/data_i[17] ,
         \words[11]/data_i[16] , \words[11]/data_i[15] ,
         \words[11]/data_i[14] , \words[11]/data_i[13] ,
         \words[11]/data_i[12] , \words[11]/data_i[11] ,
         \words[11]/data_i[10] , \words[11]/data_i[9] , \words[11]/data_i[8] ,
         \words[11]/data_i[7] , \words[11]/data_i[6] , \words[11]/data_i[5] ,
         \words[11]/data_i[4] , \words[11]/data_i[3] , \words[11]/data_i[2] ,
         \words[11]/data_i[1] , \words[11]/data_i[0] , \words[12]/valid_o ,
         \words[12]/valid_i , \words[12]/data_i[31] , \words[12]/data_i[30] ,
         \words[12]/data_i[29] , \words[12]/data_i[28] ,
         \words[12]/data_i[27] , \words[12]/data_i[26] ,
         \words[12]/data_i[25] , \words[12]/data_i[24] ,
         \words[12]/data_i[23] , \words[12]/data_i[22] ,
         \words[12]/data_i[21] , \words[12]/data_i[20] ,
         \words[12]/data_i[19] , \words[12]/data_i[18] ,
         \words[12]/data_i[17] , \words[12]/data_i[16] ,
         \words[12]/data_i[15] , \words[12]/data_i[14] ,
         \words[12]/data_i[13] , \words[12]/data_i[12] ,
         \words[12]/data_i[11] , \words[12]/data_i[10] , \words[12]/data_i[9] ,
         \words[12]/data_i[8] , \words[12]/data_i[7] , \words[12]/data_i[6] ,
         \words[12]/data_i[5] , \words[12]/data_i[4] , \words[12]/data_i[3] ,
         \words[12]/data_i[2] , \words[12]/data_i[1] , \words[12]/data_i[0] ,
         \words[13]/valid_o , \words[13]/valid_i , \words[13]/data_i[31] ,
         \words[13]/data_i[30] , \words[13]/data_i[29] ,
         \words[13]/data_i[28] , \words[13]/data_i[27] ,
         \words[13]/data_i[26] , \words[13]/data_i[25] ,
         \words[13]/data_i[24] , \words[13]/data_i[23] ,
         \words[13]/data_i[22] , \words[13]/data_i[21] ,
         \words[13]/data_i[20] , \words[13]/data_i[19] ,
         \words[13]/data_i[18] , \words[13]/data_i[17] ,
         \words[13]/data_i[16] , \words[13]/data_i[15] ,
         \words[13]/data_i[14] , \words[13]/data_i[13] ,
         \words[13]/data_i[12] , \words[13]/data_i[11] ,
         \words[13]/data_i[10] , \words[13]/data_i[9] , \words[13]/data_i[8] ,
         \words[13]/data_i[7] , \words[13]/data_i[6] , \words[13]/data_i[5] ,
         \words[13]/data_i[4] , \words[13]/data_i[3] , \words[13]/data_i[2] ,
         \words[13]/data_i[1] , \words[13]/data_i[0] , \words[14]/valid_o ,
         \words[14]/valid_i , \words[14]/data_i[31] , \words[14]/data_i[30] ,
         \words[14]/data_i[29] , \words[14]/data_i[28] ,
         \words[14]/data_i[27] , \words[14]/data_i[26] ,
         \words[14]/data_i[25] , \words[14]/data_i[24] ,
         \words[14]/data_i[23] , \words[14]/data_i[22] ,
         \words[14]/data_i[21] , \words[14]/data_i[20] ,
         \words[14]/data_i[19] , \words[14]/data_i[18] ,
         \words[14]/data_i[17] , \words[14]/data_i[16] ,
         \words[14]/data_i[15] , \words[14]/data_i[14] ,
         \words[14]/data_i[13] , \words[14]/data_i[12] ,
         \words[14]/data_i[11] , \words[14]/data_i[10] , \words[14]/data_i[9] ,
         \words[14]/data_i[8] , \words[14]/data_i[7] , \words[14]/data_i[6] ,
         \words[14]/data_i[5] , \words[14]/data_i[4] , \words[14]/data_i[3] ,
         \words[14]/data_i[2] , \words[14]/data_i[1] , \words[14]/data_i[0] ,
         \words[15]/valid_o , \words[15]/valid_i , \words[15]/data_i[31] ,
         \words[15]/data_i[30] , \words[15]/data_i[29] ,
         \words[15]/data_i[28] , \words[15]/data_i[27] ,
         \words[15]/data_i[26] , \words[15]/data_i[25] ,
         \words[15]/data_i[24] , \words[15]/data_i[23] ,
         \words[15]/data_i[22] , \words[15]/data_i[21] ,
         \words[15]/data_i[20] , \words[15]/data_i[19] ,
         \words[15]/data_i[18] , \words[15]/data_i[17] ,
         \words[15]/data_i[16] , \words[15]/data_i[15] ,
         \words[15]/data_i[14] , \words[15]/data_i[13] ,
         \words[15]/data_i[12] , \words[15]/data_i[11] ,
         \words[15]/data_i[10] , \words[15]/data_i[9] , \words[15]/data_i[8] ,
         \words[15]/data_i[7] , \words[15]/data_i[6] , \words[15]/data_i[5] ,
         \words[15]/data_i[4] , \words[15]/data_i[3] , \words[15]/data_i[2] ,
         \words[15]/data_i[1] , \words[15]/data_i[0] , \words[16]/valid_o ,
         \words[16]/valid_i , \words[16]/data_i[31] , \words[16]/data_i[30] ,
         \words[16]/data_i[29] , \words[16]/data_i[28] ,
         \words[16]/data_i[27] , \words[16]/data_i[26] ,
         \words[16]/data_i[25] , \words[16]/data_i[24] ,
         \words[16]/data_i[23] , \words[16]/data_i[22] ,
         \words[16]/data_i[21] , \words[16]/data_i[20] ,
         \words[16]/data_i[19] , \words[16]/data_i[18] ,
         \words[16]/data_i[17] , \words[16]/data_i[16] ,
         \words[16]/data_i[15] , \words[16]/data_i[14] ,
         \words[16]/data_i[13] , \words[16]/data_i[12] ,
         \words[16]/data_i[11] , \words[16]/data_i[10] , \words[16]/data_i[9] ,
         \words[16]/data_i[8] , \words[16]/data_i[7] , \words[16]/data_i[6] ,
         \words[16]/data_i[5] , \words[16]/data_i[4] , \words[16]/data_i[3] ,
         \words[16]/data_i[2] , \words[16]/data_i[1] , \words[16]/data_i[0] ,
         \words[17]/valid_o , \words[17]/valid_i , \words[17]/data_i[31] ,
         \words[17]/data_i[30] , \words[17]/data_i[29] ,
         \words[17]/data_i[28] , \words[17]/data_i[27] ,
         \words[17]/data_i[26] , \words[17]/data_i[25] ,
         \words[17]/data_i[24] , \words[17]/data_i[23] ,
         \words[17]/data_i[22] , \words[17]/data_i[21] ,
         \words[17]/data_i[20] , \words[17]/data_i[19] ,
         \words[17]/data_i[18] , \words[17]/data_i[17] ,
         \words[17]/data_i[16] , \words[17]/data_i[15] ,
         \words[17]/data_i[14] , \words[17]/data_i[13] ,
         \words[17]/data_i[12] , \words[17]/data_i[11] ,
         \words[17]/data_i[10] , \words[17]/data_i[9] , \words[17]/data_i[8] ,
         \words[17]/data_i[7] , \words[17]/data_i[6] , \words[17]/data_i[5] ,
         \words[17]/data_i[4] , \words[17]/data_i[3] , \words[17]/data_i[2] ,
         \words[17]/data_i[1] , \words[17]/data_i[0] , \words[18]/valid_o ,
         \words[18]/valid_i , \words[18]/data_i[31] , \words[18]/data_i[30] ,
         \words[18]/data_i[29] , \words[18]/data_i[28] ,
         \words[18]/data_i[27] , \words[18]/data_i[26] ,
         \words[18]/data_i[25] , \words[18]/data_i[24] ,
         \words[18]/data_i[23] , \words[18]/data_i[22] ,
         \words[18]/data_i[21] , \words[18]/data_i[20] ,
         \words[18]/data_i[19] , \words[18]/data_i[18] ,
         \words[18]/data_i[17] , \words[18]/data_i[16] ,
         \words[18]/data_i[15] , \words[18]/data_i[14] ,
         \words[18]/data_i[13] , \words[18]/data_i[12] ,
         \words[18]/data_i[11] , \words[18]/data_i[10] , \words[18]/data_i[9] ,
         \words[18]/data_i[8] , \words[18]/data_i[7] , \words[18]/data_i[6] ,
         \words[18]/data_i[5] , \words[18]/data_i[4] , \words[18]/data_i[3] ,
         \words[18]/data_i[2] , \words[18]/data_i[1] , \words[18]/data_i[0] ,
         \words[19]/valid_o , \words[19]/valid_i , \words[19]/data_i[31] ,
         \words[19]/data_i[30] , \words[19]/data_i[29] ,
         \words[19]/data_i[28] , \words[19]/data_i[27] ,
         \words[19]/data_i[26] , \words[19]/data_i[25] ,
         \words[19]/data_i[24] , \words[19]/data_i[23] ,
         \words[19]/data_i[22] , \words[19]/data_i[21] ,
         \words[19]/data_i[20] , \words[19]/data_i[19] ,
         \words[19]/data_i[18] , \words[19]/data_i[17] ,
         \words[19]/data_i[16] , \words[19]/data_i[15] ,
         \words[19]/data_i[14] , \words[19]/data_i[13] ,
         \words[19]/data_i[12] , \words[19]/data_i[11] ,
         \words[19]/data_i[10] , \words[19]/data_i[9] , \words[19]/data_i[8] ,
         \words[19]/data_i[7] , \words[19]/data_i[6] , \words[19]/data_i[5] ,
         \words[19]/data_i[4] , \words[19]/data_i[3] , \words[19]/data_i[2] ,
         \words[19]/data_i[1] , \words[19]/data_i[0] , \words[20]/valid_o ,
         \words[20]/valid_i , \words[20]/data_i[31] , \words[20]/data_i[30] ,
         \words[20]/data_i[29] , \words[20]/data_i[28] ,
         \words[20]/data_i[27] , \words[20]/data_i[26] ,
         \words[20]/data_i[25] , \words[20]/data_i[24] ,
         \words[20]/data_i[23] , \words[20]/data_i[22] ,
         \words[20]/data_i[21] , \words[20]/data_i[20] ,
         \words[20]/data_i[19] , \words[20]/data_i[18] ,
         \words[20]/data_i[17] , \words[20]/data_i[16] ,
         \words[20]/data_i[15] , \words[20]/data_i[14] ,
         \words[20]/data_i[13] , \words[20]/data_i[12] ,
         \words[20]/data_i[11] , \words[20]/data_i[10] , \words[20]/data_i[9] ,
         \words[20]/data_i[8] , \words[20]/data_i[7] , \words[20]/data_i[6] ,
         \words[20]/data_i[5] , \words[20]/data_i[4] , \words[20]/data_i[3] ,
         \words[20]/data_i[2] , \words[20]/data_i[1] , \words[20]/data_i[0] ,
         \words[21]/valid_o , \words[21]/valid_i , \words[21]/data_i[31] ,
         \words[21]/data_i[30] , \words[21]/data_i[29] ,
         \words[21]/data_i[28] , \words[21]/data_i[27] ,
         \words[21]/data_i[26] , \words[21]/data_i[25] ,
         \words[21]/data_i[24] , \words[21]/data_i[23] ,
         \words[21]/data_i[22] , \words[21]/data_i[21] ,
         \words[21]/data_i[20] , \words[21]/data_i[19] ,
         \words[21]/data_i[18] , \words[21]/data_i[17] ,
         \words[21]/data_i[16] , \words[21]/data_i[15] ,
         \words[21]/data_i[14] , \words[21]/data_i[13] ,
         \words[21]/data_i[12] , \words[21]/data_i[11] ,
         \words[21]/data_i[10] , \words[21]/data_i[9] , \words[21]/data_i[8] ,
         \words[21]/data_i[7] , \words[21]/data_i[6] , \words[21]/data_i[5] ,
         \words[21]/data_i[4] , \words[21]/data_i[3] , \words[21]/data_i[2] ,
         \words[21]/data_i[1] , \words[21]/data_i[0] , \words[22]/valid_o ,
         \words[22]/valid_i , \words[22]/data_i[31] , \words[22]/data_i[30] ,
         \words[22]/data_i[29] , \words[22]/data_i[28] ,
         \words[22]/data_i[27] , \words[22]/data_i[26] ,
         \words[22]/data_i[25] , \words[22]/data_i[24] ,
         \words[22]/data_i[23] , \words[22]/data_i[22] ,
         \words[22]/data_i[21] , \words[22]/data_i[20] ,
         \words[22]/data_i[19] , \words[22]/data_i[18] ,
         \words[22]/data_i[17] , \words[22]/data_i[16] ,
         \words[22]/data_i[15] , \words[22]/data_i[14] ,
         \words[22]/data_i[13] , \words[22]/data_i[12] ,
         \words[22]/data_i[11] , \words[22]/data_i[10] , \words[22]/data_i[9] ,
         \words[22]/data_i[8] , \words[22]/data_i[7] , \words[22]/data_i[6] ,
         \words[22]/data_i[5] , \words[22]/data_i[4] , \words[22]/data_i[3] ,
         \words[22]/data_i[2] , \words[22]/data_i[1] , \words[22]/data_i[0] ,
         \words[23]/valid_o , \words[23]/valid_i , \words[23]/data_i[31] ,
         \words[23]/data_i[30] , \words[23]/data_i[29] ,
         \words[23]/data_i[28] , \words[23]/data_i[27] ,
         \words[23]/data_i[26] , \words[23]/data_i[25] ,
         \words[23]/data_i[24] , \words[23]/data_i[23] ,
         \words[23]/data_i[22] , \words[23]/data_i[21] ,
         \words[23]/data_i[20] , \words[23]/data_i[19] ,
         \words[23]/data_i[18] , \words[23]/data_i[17] ,
         \words[23]/data_i[16] , \words[23]/data_i[15] ,
         \words[23]/data_i[14] , \words[23]/data_i[13] ,
         \words[23]/data_i[12] , \words[23]/data_i[11] ,
         \words[23]/data_i[10] , \words[23]/data_i[9] , \words[23]/data_i[8] ,
         \words[23]/data_i[7] , \words[23]/data_i[6] , \words[23]/data_i[5] ,
         \words[23]/data_i[4] , \words[23]/data_i[3] , \words[23]/data_i[2] ,
         \words[23]/data_i[1] , \words[23]/data_i[0] , \words[24]/valid_o ,
         \words[24]/valid_i , \words[24]/data_i[31] , \words[24]/data_i[30] ,
         \words[24]/data_i[29] , \words[24]/data_i[28] ,
         \words[24]/data_i[27] , \words[24]/data_i[26] ,
         \words[24]/data_i[25] , \words[24]/data_i[24] ,
         \words[24]/data_i[23] , \words[24]/data_i[22] ,
         \words[24]/data_i[21] , \words[24]/data_i[20] ,
         \words[24]/data_i[19] , \words[24]/data_i[18] ,
         \words[24]/data_i[17] , \words[24]/data_i[16] ,
         \words[24]/data_i[15] , \words[24]/data_i[14] ,
         \words[24]/data_i[13] , \words[24]/data_i[12] ,
         \words[24]/data_i[11] , \words[24]/data_i[10] , \words[24]/data_i[9] ,
         \words[24]/data_i[8] , \words[24]/data_i[7] , \words[24]/data_i[6] ,
         \words[24]/data_i[5] , \words[24]/data_i[4] , \words[24]/data_i[3] ,
         \words[24]/data_i[2] , \words[24]/data_i[1] , \words[24]/data_i[0] ,
         \words[25]/valid_o , \words[25]/valid_i , \words[25]/data_i[31] ,
         \words[25]/data_i[30] , \words[25]/data_i[29] ,
         \words[25]/data_i[28] , \words[25]/data_i[27] ,
         \words[25]/data_i[26] , \words[25]/data_i[25] ,
         \words[25]/data_i[24] , \words[25]/data_i[23] ,
         \words[25]/data_i[22] , \words[25]/data_i[21] ,
         \words[25]/data_i[20] , \words[25]/data_i[19] ,
         \words[25]/data_i[18] , \words[25]/data_i[17] ,
         \words[25]/data_i[16] , \words[25]/data_i[15] ,
         \words[25]/data_i[14] , \words[25]/data_i[13] ,
         \words[25]/data_i[12] , \words[25]/data_i[11] ,
         \words[25]/data_i[10] , \words[25]/data_i[9] , \words[25]/data_i[8] ,
         \words[25]/data_i[7] , \words[25]/data_i[6] , \words[25]/data_i[5] ,
         \words[25]/data_i[4] , \words[25]/data_i[3] , \words[25]/data_i[2] ,
         \words[25]/data_i[1] , \words[25]/data_i[0] , \words[26]/valid_o ,
         \words[26]/valid_i , \words[26]/data_i[31] , \words[26]/data_i[30] ,
         \words[26]/data_i[29] , \words[26]/data_i[28] ,
         \words[26]/data_i[27] , \words[26]/data_i[26] ,
         \words[26]/data_i[25] , \words[26]/data_i[24] ,
         \words[26]/data_i[23] , \words[26]/data_i[22] ,
         \words[26]/data_i[21] , \words[26]/data_i[20] ,
         \words[26]/data_i[19] , \words[26]/data_i[18] ,
         \words[26]/data_i[17] , \words[26]/data_i[16] ,
         \words[26]/data_i[15] , \words[26]/data_i[14] ,
         \words[26]/data_i[13] , \words[26]/data_i[12] ,
         \words[26]/data_i[11] , \words[26]/data_i[10] , \words[26]/data_i[9] ,
         \words[26]/data_i[8] , \words[26]/data_i[7] , \words[26]/data_i[6] ,
         \words[26]/data_i[5] , \words[26]/data_i[4] , \words[26]/data_i[3] ,
         \words[26]/data_i[2] , \words[26]/data_i[1] , \words[26]/data_i[0] ,
         \words[27]/valid_o , \words[27]/valid_i , \words[27]/data_i[31] ,
         \words[27]/data_i[30] , \words[27]/data_i[29] ,
         \words[27]/data_i[28] , \words[27]/data_i[27] ,
         \words[27]/data_i[26] , \words[27]/data_i[25] ,
         \words[27]/data_i[24] , \words[27]/data_i[23] ,
         \words[27]/data_i[22] , \words[27]/data_i[21] ,
         \words[27]/data_i[20] , \words[27]/data_i[19] ,
         \words[27]/data_i[18] , \words[27]/data_i[17] ,
         \words[27]/data_i[16] , \words[27]/data_i[15] ,
         \words[27]/data_i[14] , \words[27]/data_i[13] ,
         \words[27]/data_i[12] , \words[27]/data_i[11] ,
         \words[27]/data_i[10] , \words[27]/data_i[9] , \words[27]/data_i[8] ,
         \words[27]/data_i[7] , \words[27]/data_i[6] , \words[27]/data_i[5] ,
         \words[27]/data_i[4] , \words[27]/data_i[3] , \words[27]/data_i[2] ,
         \words[27]/data_i[1] , \words[27]/data_i[0] , \words[28]/valid_o ,
         \words[28]/valid_i , \words[28]/data_i[31] , \words[28]/data_i[30] ,
         \words[28]/data_i[29] , \words[28]/data_i[28] ,
         \words[28]/data_i[27] , \words[28]/data_i[26] ,
         \words[28]/data_i[25] , \words[28]/data_i[24] ,
         \words[28]/data_i[23] , \words[28]/data_i[22] ,
         \words[28]/data_i[21] , \words[28]/data_i[20] ,
         \words[28]/data_i[19] , \words[28]/data_i[18] ,
         \words[28]/data_i[17] , \words[28]/data_i[16] ,
         \words[28]/data_i[15] , \words[28]/data_i[14] ,
         \words[28]/data_i[13] , \words[28]/data_i[12] ,
         \words[28]/data_i[11] , \words[28]/data_i[10] , \words[28]/data_i[9] ,
         \words[28]/data_i[8] , \words[28]/data_i[7] , \words[28]/data_i[6] ,
         \words[28]/data_i[5] , \words[28]/data_i[4] , \words[28]/data_i[3] ,
         \words[28]/data_i[2] , \words[28]/data_i[1] , \words[28]/data_i[0] ,
         \words[29]/valid_o , \words[29]/valid_i , \words[29]/data_i[31] ,
         \words[29]/data_i[30] , \words[29]/data_i[29] ,
         \words[29]/data_i[28] , \words[29]/data_i[27] ,
         \words[29]/data_i[26] , \words[29]/data_i[25] ,
         \words[29]/data_i[24] , \words[29]/data_i[23] ,
         \words[29]/data_i[22] , \words[29]/data_i[21] ,
         \words[29]/data_i[20] , \words[29]/data_i[19] ,
         \words[29]/data_i[18] , \words[29]/data_i[17] ,
         \words[29]/data_i[16] , \words[29]/data_i[15] ,
         \words[29]/data_i[14] , \words[29]/data_i[13] ,
         \words[29]/data_i[12] , \words[29]/data_i[11] ,
         \words[29]/data_i[10] , \words[29]/data_i[9] , \words[29]/data_i[8] ,
         \words[29]/data_i[7] , \words[29]/data_i[6] , \words[29]/data_i[5] ,
         \words[29]/data_i[4] , \words[29]/data_i[3] , \words[29]/data_i[2] ,
         \words[29]/data_i[1] , \words[29]/data_i[0] , \words[30]/valid_o ,
         \words[30]/valid_i , \words[30]/data_i[31] , \words[30]/data_i[30] ,
         \words[30]/data_i[29] , \words[30]/data_i[28] ,
         \words[30]/data_i[27] , \words[30]/data_i[26] ,
         \words[30]/data_i[25] , \words[30]/data_i[24] ,
         \words[30]/data_i[23] , \words[30]/data_i[22] ,
         \words[30]/data_i[21] , \words[30]/data_i[20] ,
         \words[30]/data_i[19] , \words[30]/data_i[18] ,
         \words[30]/data_i[17] , \words[30]/data_i[16] ,
         \words[30]/data_i[15] , \words[30]/data_i[14] ,
         \words[30]/data_i[13] , \words[30]/data_i[12] ,
         \words[30]/data_i[11] , \words[30]/data_i[10] , \words[30]/data_i[9] ,
         \words[30]/data_i[8] , \words[30]/data_i[7] , \words[30]/data_i[6] ,
         \words[30]/data_i[5] , \words[30]/data_i[4] , \words[30]/data_i[3] ,
         \words[30]/data_i[2] , \words[30]/data_i[1] , \words[30]/data_i[0] ,
         n6, n7, n11, n12, n14, n15, n16, n17, n18, n19, n21, n22, n23, n24,
         n26, n27, n28, n29, n30, n31, n34, n37, n38, n39, n40, n43, n44, n45,
         n46, n48, n49, n50, n51, n53, n54, n55, n56, n58, n59, n60, n61, n64,
         n65, n66, n67, n69, n70, n71, n72, n74, n75, n76, n77, n79, n80, n81,
         n82, n83, n84, n85, n86, n88, n89, n1480, n1481, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1494, n1495, n1496,
         n1497, n1498, n1499, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115;

  mux read_mux ( .data_i({\read_value_mux[31][31] , \read_value_mux[31][30] , 
        \read_value_mux[31][29] , \read_value_mux[31][28] , 
        \read_value_mux[31][27] , \read_value_mux[31][26] , 
        \read_value_mux[31][25] , \read_value_mux[31][24] , 
        \read_value_mux[31][23] , \read_value_mux[31][22] , 
        \read_value_mux[31][21] , \read_value_mux[31][20] , 
        \read_value_mux[31][19] , \read_value_mux[31][18] , 
        \read_value_mux[31][17] , \read_value_mux[31][16] , 
        \read_value_mux[31][15] , \read_value_mux[31][14] , 
        \read_value_mux[31][13] , \read_value_mux[31][12] , 
        \read_value_mux[31][11] , \read_value_mux[31][10] , 
        \read_value_mux[31][9] , \read_value_mux[31][8] , 
        \read_value_mux[31][7] , \read_value_mux[31][6] , 
        \read_value_mux[31][5] , \read_value_mux[31][4] , 
        \read_value_mux[31][3] , \read_value_mux[31][2] , 
        \read_value_mux[31][1] , \read_value_mux[31][0] , 
        \read_value_mux[30][31] , \read_value_mux[30][30] , 
        \read_value_mux[30][29] , \read_value_mux[30][28] , 
        \read_value_mux[30][27] , \read_value_mux[30][26] , 
        \read_value_mux[30][25] , \read_value_mux[30][24] , 
        \read_value_mux[30][23] , \read_value_mux[30][22] , 
        \read_value_mux[30][21] , \read_value_mux[30][20] , 
        \read_value_mux[30][19] , \read_value_mux[30][18] , 
        \read_value_mux[30][17] , \read_value_mux[30][16] , 
        \read_value_mux[30][15] , \read_value_mux[30][14] , 
        \read_value_mux[30][13] , \read_value_mux[30][12] , 
        \read_value_mux[30][11] , \read_value_mux[30][10] , 
        \read_value_mux[30][9] , \read_value_mux[30][8] , 
        \read_value_mux[30][7] , \read_value_mux[30][6] , 
        \read_value_mux[30][5] , \read_value_mux[30][4] , 
        \read_value_mux[30][3] , \read_value_mux[30][2] , 
        \read_value_mux[30][1] , \read_value_mux[30][0] , 
        \read_value_mux[29][31] , \read_value_mux[29][30] , 
        \read_value_mux[29][29] , \read_value_mux[29][28] , 
        \read_value_mux[29][27] , \read_value_mux[29][26] , 
        \read_value_mux[29][25] , \read_value_mux[29][24] , 
        \read_value_mux[29][23] , \read_value_mux[29][22] , 
        \read_value_mux[29][21] , \read_value_mux[29][20] , 
        \read_value_mux[29][19] , \read_value_mux[29][18] , 
        \read_value_mux[29][17] , \read_value_mux[29][16] , 
        \read_value_mux[29][15] , \read_value_mux[29][14] , 
        \read_value_mux[29][13] , \read_value_mux[29][12] , 
        \read_value_mux[29][11] , \read_value_mux[29][10] , 
        \read_value_mux[29][9] , \read_value_mux[29][8] , 
        \read_value_mux[29][7] , \read_value_mux[29][6] , 
        \read_value_mux[29][5] , \read_value_mux[29][4] , 
        \read_value_mux[29][3] , \read_value_mux[29][2] , 
        \read_value_mux[29][1] , \read_value_mux[29][0] , 
        \read_value_mux[28][31] , \read_value_mux[28][30] , 
        \read_value_mux[28][29] , \read_value_mux[28][28] , 
        \read_value_mux[28][27] , \read_value_mux[28][26] , 
        \read_value_mux[28][25] , \read_value_mux[28][24] , 
        \read_value_mux[28][23] , \read_value_mux[28][22] , 
        \read_value_mux[28][21] , \read_value_mux[28][20] , 
        \read_value_mux[28][19] , \read_value_mux[28][18] , 
        \read_value_mux[28][17] , \read_value_mux[28][16] , 
        \read_value_mux[28][15] , \read_value_mux[28][14] , 
        \read_value_mux[28][13] , \read_value_mux[28][12] , 
        \read_value_mux[28][11] , \read_value_mux[28][10] , 
        \read_value_mux[28][9] , \read_value_mux[28][8] , 
        \read_value_mux[28][7] , \read_value_mux[28][6] , 
        \read_value_mux[28][5] , \read_value_mux[28][4] , 
        \read_value_mux[28][3] , \read_value_mux[28][2] , 
        \read_value_mux[28][1] , \read_value_mux[28][0] , 
        \read_value_mux[27][31] , \read_value_mux[27][30] , 
        \read_value_mux[27][29] , \read_value_mux[27][28] , 
        \read_value_mux[27][27] , \read_value_mux[27][26] , 
        \read_value_mux[27][25] , \read_value_mux[27][24] , 
        \read_value_mux[27][23] , \read_value_mux[27][22] , 
        \read_value_mux[27][21] , \read_value_mux[27][20] , 
        \read_value_mux[27][19] , \read_value_mux[27][18] , 
        \read_value_mux[27][17] , \read_value_mux[27][16] , 
        \read_value_mux[27][15] , \read_value_mux[27][14] , 
        \read_value_mux[27][13] , \read_value_mux[27][12] , 
        \read_value_mux[27][11] , \read_value_mux[27][10] , 
        \read_value_mux[27][9] , \read_value_mux[27][8] , 
        \read_value_mux[27][7] , \read_value_mux[27][6] , 
        \read_value_mux[27][5] , \read_value_mux[27][4] , 
        \read_value_mux[27][3] , \read_value_mux[27][2] , 
        \read_value_mux[27][1] , \read_value_mux[27][0] , 
        \read_value_mux[26][31] , \read_value_mux[26][30] , 
        \read_value_mux[26][29] , \read_value_mux[26][28] , 
        \read_value_mux[26][27] , \read_value_mux[26][26] , 
        \read_value_mux[26][25] , \read_value_mux[26][24] , 
        \read_value_mux[26][23] , \read_value_mux[26][22] , 
        \read_value_mux[26][21] , \read_value_mux[26][20] , 
        \read_value_mux[26][19] , \read_value_mux[26][18] , 
        \read_value_mux[26][17] , \read_value_mux[26][16] , 
        \read_value_mux[26][15] , \read_value_mux[26][14] , 
        \read_value_mux[26][13] , \read_value_mux[26][12] , 
        \read_value_mux[26][11] , \read_value_mux[26][10] , 
        \read_value_mux[26][9] , \read_value_mux[26][8] , 
        \read_value_mux[26][7] , \read_value_mux[26][6] , 
        \read_value_mux[26][5] , \read_value_mux[26][4] , 
        \read_value_mux[26][3] , \read_value_mux[26][2] , 
        \read_value_mux[26][1] , \read_value_mux[26][0] , 
        \read_value_mux[25][31] , \read_value_mux[25][30] , 
        \read_value_mux[25][29] , \read_value_mux[25][28] , 
        \read_value_mux[25][27] , \read_value_mux[25][26] , 
        \read_value_mux[25][25] , \read_value_mux[25][24] , 
        \read_value_mux[25][23] , \read_value_mux[25][22] , 
        \read_value_mux[25][21] , \read_value_mux[25][20] , 
        \read_value_mux[25][19] , \read_value_mux[25][18] , 
        \read_value_mux[25][17] , \read_value_mux[25][16] , 
        \read_value_mux[25][15] , \read_value_mux[25][14] , 
        \read_value_mux[25][13] , \read_value_mux[25][12] , 
        \read_value_mux[25][11] , \read_value_mux[25][10] , 
        \read_value_mux[25][9] , \read_value_mux[25][8] , 
        \read_value_mux[25][7] , \read_value_mux[25][6] , 
        \read_value_mux[25][5] , \read_value_mux[25][4] , 
        \read_value_mux[25][3] , \read_value_mux[25][2] , 
        \read_value_mux[25][1] , \read_value_mux[25][0] , 
        \read_value_mux[24][31] , \read_value_mux[24][30] , 
        \read_value_mux[24][29] , \read_value_mux[24][28] , 
        \read_value_mux[24][27] , \read_value_mux[24][26] , 
        \read_value_mux[24][25] , \read_value_mux[24][24] , 
        \read_value_mux[24][23] , \read_value_mux[24][22] , 
        \read_value_mux[24][21] , \read_value_mux[24][20] , 
        \read_value_mux[24][19] , \read_value_mux[24][18] , 
        \read_value_mux[24][17] , \read_value_mux[24][16] , 
        \read_value_mux[24][15] , \read_value_mux[24][14] , 
        \read_value_mux[24][13] , \read_value_mux[24][12] , 
        \read_value_mux[24][11] , \read_value_mux[24][10] , 
        \read_value_mux[24][9] , \read_value_mux[24][8] , 
        \read_value_mux[24][7] , \read_value_mux[24][6] , 
        \read_value_mux[24][5] , \read_value_mux[24][4] , 
        \read_value_mux[24][3] , \read_value_mux[24][2] , 
        \read_value_mux[24][1] , \read_value_mux[24][0] , 
        \read_value_mux[23][31] , \read_value_mux[23][30] , 
        \read_value_mux[23][29] , \read_value_mux[23][28] , 
        \read_value_mux[23][27] , \read_value_mux[23][26] , 
        \read_value_mux[23][25] , \read_value_mux[23][24] , 
        \read_value_mux[23][23] , \read_value_mux[23][22] , 
        \read_value_mux[23][21] , \read_value_mux[23][20] , 
        \read_value_mux[23][19] , \read_value_mux[23][18] , 
        \read_value_mux[23][17] , \read_value_mux[23][16] , 
        \read_value_mux[23][15] , \read_value_mux[23][14] , 
        \read_value_mux[23][13] , \read_value_mux[23][12] , 
        \read_value_mux[23][11] , \read_value_mux[23][10] , 
        \read_value_mux[23][9] , \read_value_mux[23][8] , 
        \read_value_mux[23][7] , \read_value_mux[23][6] , 
        \read_value_mux[23][5] , \read_value_mux[23][4] , 
        \read_value_mux[23][3] , \read_value_mux[23][2] , 
        \read_value_mux[23][1] , \read_value_mux[23][0] , 
        \read_value_mux[22][31] , \read_value_mux[22][30] , 
        \read_value_mux[22][29] , \read_value_mux[22][28] , 
        \read_value_mux[22][27] , \read_value_mux[22][26] , 
        \read_value_mux[22][25] , \read_value_mux[22][24] , 
        \read_value_mux[22][23] , \read_value_mux[22][22] , 
        \read_value_mux[22][21] , \read_value_mux[22][20] , 
        \read_value_mux[22][19] , \read_value_mux[22][18] , 
        \read_value_mux[22][17] , \read_value_mux[22][16] , 
        \read_value_mux[22][15] , \read_value_mux[22][14] , 
        \read_value_mux[22][13] , \read_value_mux[22][12] , 
        \read_value_mux[22][11] , \read_value_mux[22][10] , 
        \read_value_mux[22][9] , \read_value_mux[22][8] , 
        \read_value_mux[22][7] , \read_value_mux[22][6] , 
        \read_value_mux[22][5] , \read_value_mux[22][4] , 
        \read_value_mux[22][3] , \read_value_mux[22][2] , 
        \read_value_mux[22][1] , \read_value_mux[22][0] , 
        \read_value_mux[21][31] , \read_value_mux[21][30] , 
        \read_value_mux[21][29] , \read_value_mux[21][28] , 
        \read_value_mux[21][27] , \read_value_mux[21][26] , 
        \read_value_mux[21][25] , \read_value_mux[21][24] , 
        \read_value_mux[21][23] , \read_value_mux[21][22] , 
        \read_value_mux[21][21] , \read_value_mux[21][20] , 
        \read_value_mux[21][19] , \read_value_mux[21][18] , 
        \read_value_mux[21][17] , \read_value_mux[21][16] , 
        \read_value_mux[21][15] , \read_value_mux[21][14] , 
        \read_value_mux[21][13] , \read_value_mux[21][12] , 
        \read_value_mux[21][11] , \read_value_mux[21][10] , 
        \read_value_mux[21][9] , \read_value_mux[21][8] , 
        \read_value_mux[21][7] , \read_value_mux[21][6] , 
        \read_value_mux[21][5] , \read_value_mux[21][4] , 
        \read_value_mux[21][3] , \read_value_mux[21][2] , 
        \read_value_mux[21][1] , \read_value_mux[21][0] , 
        \read_value_mux[20][31] , \read_value_mux[20][30] , 
        \read_value_mux[20][29] , \read_value_mux[20][28] , 
        \read_value_mux[20][27] , \read_value_mux[20][26] , 
        \read_value_mux[20][25] , \read_value_mux[20][24] , 
        \read_value_mux[20][23] , \read_value_mux[20][22] , 
        \read_value_mux[20][21] , \read_value_mux[20][20] , 
        \read_value_mux[20][19] , \read_value_mux[20][18] , 
        \read_value_mux[20][17] , \read_value_mux[20][16] , 
        \read_value_mux[20][15] , \read_value_mux[20][14] , 
        \read_value_mux[20][13] , \read_value_mux[20][12] , 
        \read_value_mux[20][11] , \read_value_mux[20][10] , 
        \read_value_mux[20][9] , \read_value_mux[20][8] , 
        \read_value_mux[20][7] , \read_value_mux[20][6] , 
        \read_value_mux[20][5] , \read_value_mux[20][4] , 
        \read_value_mux[20][3] , \read_value_mux[20][2] , 
        \read_value_mux[20][1] , \read_value_mux[20][0] , 
        \read_value_mux[19][31] , \read_value_mux[19][30] , 
        \read_value_mux[19][29] , \read_value_mux[19][28] , 
        \read_value_mux[19][27] , \read_value_mux[19][26] , 
        \read_value_mux[19][25] , \read_value_mux[19][24] , 
        \read_value_mux[19][23] , \read_value_mux[19][22] , 
        \read_value_mux[19][21] , \read_value_mux[19][20] , 
        \read_value_mux[19][19] , \read_value_mux[19][18] , 
        \read_value_mux[19][17] , \read_value_mux[19][16] , 
        \read_value_mux[19][15] , \read_value_mux[19][14] , 
        \read_value_mux[19][13] , \read_value_mux[19][12] , 
        \read_value_mux[19][11] , \read_value_mux[19][10] , 
        \read_value_mux[19][9] , \read_value_mux[19][8] , 
        \read_value_mux[19][7] , \read_value_mux[19][6] , 
        \read_value_mux[19][5] , \read_value_mux[19][4] , 
        \read_value_mux[19][3] , \read_value_mux[19][2] , 
        \read_value_mux[19][1] , \read_value_mux[19][0] , 
        \read_value_mux[18][31] , \read_value_mux[18][30] , 
        \read_value_mux[18][29] , \read_value_mux[18][28] , 
        \read_value_mux[18][27] , \read_value_mux[18][26] , 
        \read_value_mux[18][25] , \read_value_mux[18][24] , 
        \read_value_mux[18][23] , \read_value_mux[18][22] , 
        \read_value_mux[18][21] , \read_value_mux[18][20] , 
        \read_value_mux[18][19] , \read_value_mux[18][18] , 
        \read_value_mux[18][17] , \read_value_mux[18][16] , 
        \read_value_mux[18][15] , \read_value_mux[18][14] , 
        \read_value_mux[18][13] , \read_value_mux[18][12] , 
        \read_value_mux[18][11] , \read_value_mux[18][10] , 
        \read_value_mux[18][9] , \read_value_mux[18][8] , 
        \read_value_mux[18][7] , \read_value_mux[18][6] , 
        \read_value_mux[18][5] , \read_value_mux[18][4] , 
        \read_value_mux[18][3] , \read_value_mux[18][2] , 
        \read_value_mux[18][1] , \read_value_mux[18][0] , 
        \read_value_mux[17][31] , \read_value_mux[17][30] , 
        \read_value_mux[17][29] , \read_value_mux[17][28] , 
        \read_value_mux[17][27] , \read_value_mux[17][26] , 
        \read_value_mux[17][25] , \read_value_mux[17][24] , 
        \read_value_mux[17][23] , \read_value_mux[17][22] , 
        \read_value_mux[17][21] , \read_value_mux[17][20] , 
        \read_value_mux[17][19] , \read_value_mux[17][18] , 
        \read_value_mux[17][17] , \read_value_mux[17][16] , 
        \read_value_mux[17][15] , \read_value_mux[17][14] , 
        \read_value_mux[17][13] , \read_value_mux[17][12] , 
        \read_value_mux[17][11] , \read_value_mux[17][10] , 
        \read_value_mux[17][9] , \read_value_mux[17][8] , 
        \read_value_mux[17][7] , \read_value_mux[17][6] , 
        \read_value_mux[17][5] , \read_value_mux[17][4] , 
        \read_value_mux[17][3] , \read_value_mux[17][2] , 
        \read_value_mux[17][1] , \read_value_mux[17][0] , 
        \read_value_mux[16][31] , \read_value_mux[16][30] , 
        \read_value_mux[16][29] , \read_value_mux[16][28] , 
        \read_value_mux[16][27] , \read_value_mux[16][26] , 
        \read_value_mux[16][25] , \read_value_mux[16][24] , 
        \read_value_mux[16][23] , \read_value_mux[16][22] , 
        \read_value_mux[16][21] , \read_value_mux[16][20] , 
        \read_value_mux[16][19] , \read_value_mux[16][18] , 
        \read_value_mux[16][17] , \read_value_mux[16][16] , 
        \read_value_mux[16][15] , \read_value_mux[16][14] , 
        \read_value_mux[16][13] , \read_value_mux[16][12] , 
        \read_value_mux[16][11] , \read_value_mux[16][10] , 
        \read_value_mux[16][9] , \read_value_mux[16][8] , 
        \read_value_mux[16][7] , \read_value_mux[16][6] , 
        \read_value_mux[16][5] , \read_value_mux[16][4] , 
        \read_value_mux[16][3] , \read_value_mux[16][2] , 
        \read_value_mux[16][1] , \read_value_mux[16][0] , 
        \read_value_mux[15][31] , \read_value_mux[15][30] , 
        \read_value_mux[15][29] , \read_value_mux[15][28] , 
        \read_value_mux[15][27] , \read_value_mux[15][26] , 
        \read_value_mux[15][25] , \read_value_mux[15][24] , 
        \read_value_mux[15][23] , \read_value_mux[15][22] , 
        \read_value_mux[15][21] , \read_value_mux[15][20] , 
        \read_value_mux[15][19] , \read_value_mux[15][18] , 
        \read_value_mux[15][17] , \read_value_mux[15][16] , 
        \read_value_mux[15][15] , \read_value_mux[15][14] , 
        \read_value_mux[15][13] , \read_value_mux[15][12] , 
        \read_value_mux[15][11] , \read_value_mux[15][10] , 
        \read_value_mux[15][9] , \read_value_mux[15][8] , 
        \read_value_mux[15][7] , \read_value_mux[15][6] , 
        \read_value_mux[15][5] , \read_value_mux[15][4] , 
        \read_value_mux[15][3] , \read_value_mux[15][2] , 
        \read_value_mux[15][1] , \read_value_mux[15][0] , 
        \read_value_mux[14][31] , \read_value_mux[14][30] , 
        \read_value_mux[14][29] , \read_value_mux[14][28] , 
        \read_value_mux[14][27] , \read_value_mux[14][26] , 
        \read_value_mux[14][25] , \read_value_mux[14][24] , 
        \read_value_mux[14][23] , \read_value_mux[14][22] , 
        \read_value_mux[14][21] , \read_value_mux[14][20] , 
        \read_value_mux[14][19] , \read_value_mux[14][18] , 
        \read_value_mux[14][17] , \read_value_mux[14][16] , 
        \read_value_mux[14][15] , \read_value_mux[14][14] , 
        \read_value_mux[14][13] , \read_value_mux[14][12] , 
        \read_value_mux[14][11] , \read_value_mux[14][10] , 
        \read_value_mux[14][9] , \read_value_mux[14][8] , 
        \read_value_mux[14][7] , \read_value_mux[14][6] , 
        \read_value_mux[14][5] , \read_value_mux[14][4] , 
        \read_value_mux[14][3] , \read_value_mux[14][2] , 
        \read_value_mux[14][1] , \read_value_mux[14][0] , 
        \read_value_mux[13][31] , \read_value_mux[13][30] , 
        \read_value_mux[13][29] , \read_value_mux[13][28] , 
        \read_value_mux[13][27] , \read_value_mux[13][26] , 
        \read_value_mux[13][25] , \read_value_mux[13][24] , 
        \read_value_mux[13][23] , \read_value_mux[13][22] , 
        \read_value_mux[13][21] , \read_value_mux[13][20] , 
        \read_value_mux[13][19] , \read_value_mux[13][18] , 
        \read_value_mux[13][17] , \read_value_mux[13][16] , 
        \read_value_mux[13][15] , \read_value_mux[13][14] , 
        \read_value_mux[13][13] , \read_value_mux[13][12] , 
        \read_value_mux[13][11] , \read_value_mux[13][10] , 
        \read_value_mux[13][9] , \read_value_mux[13][8] , 
        \read_value_mux[13][7] , \read_value_mux[13][6] , 
        \read_value_mux[13][5] , \read_value_mux[13][4] , 
        \read_value_mux[13][3] , \read_value_mux[13][2] , 
        \read_value_mux[13][1] , \read_value_mux[13][0] , 
        \read_value_mux[12][31] , \read_value_mux[12][30] , 
        \read_value_mux[12][29] , \read_value_mux[12][28] , 
        \read_value_mux[12][27] , \read_value_mux[12][26] , 
        \read_value_mux[12][25] , \read_value_mux[12][24] , 
        \read_value_mux[12][23] , \read_value_mux[12][22] , 
        \read_value_mux[12][21] , \read_value_mux[12][20] , 
        \read_value_mux[12][19] , \read_value_mux[12][18] , 
        \read_value_mux[12][17] , \read_value_mux[12][16] , 
        \read_value_mux[12][15] , \read_value_mux[12][14] , 
        \read_value_mux[12][13] , \read_value_mux[12][12] , 
        \read_value_mux[12][11] , \read_value_mux[12][10] , 
        \read_value_mux[12][9] , \read_value_mux[12][8] , 
        \read_value_mux[12][7] , \read_value_mux[12][6] , 
        \read_value_mux[12][5] , \read_value_mux[12][4] , 
        \read_value_mux[12][3] , \read_value_mux[12][2] , 
        \read_value_mux[12][1] , \read_value_mux[12][0] , 
        \read_value_mux[11][31] , \read_value_mux[11][30] , 
        \read_value_mux[11][29] , \read_value_mux[11][28] , 
        \read_value_mux[11][27] , \read_value_mux[11][26] , 
        \read_value_mux[11][25] , \read_value_mux[11][24] , 
        \read_value_mux[11][23] , \read_value_mux[11][22] , 
        \read_value_mux[11][21] , \read_value_mux[11][20] , 
        \read_value_mux[11][19] , \read_value_mux[11][18] , 
        \read_value_mux[11][17] , \read_value_mux[11][16] , 
        \read_value_mux[11][15] , \read_value_mux[11][14] , 
        \read_value_mux[11][13] , \read_value_mux[11][12] , 
        \read_value_mux[11][11] , \read_value_mux[11][10] , 
        \read_value_mux[11][9] , \read_value_mux[11][8] , 
        \read_value_mux[11][7] , \read_value_mux[11][6] , 
        \read_value_mux[11][5] , \read_value_mux[11][4] , 
        \read_value_mux[11][3] , \read_value_mux[11][2] , 
        \read_value_mux[11][1] , \read_value_mux[11][0] , 
        \read_value_mux[10][31] , \read_value_mux[10][30] , 
        \read_value_mux[10][29] , \read_value_mux[10][28] , 
        \read_value_mux[10][27] , \read_value_mux[10][26] , 
        \read_value_mux[10][25] , \read_value_mux[10][24] , 
        \read_value_mux[10][23] , \read_value_mux[10][22] , 
        \read_value_mux[10][21] , \read_value_mux[10][20] , 
        \read_value_mux[10][19] , \read_value_mux[10][18] , 
        \read_value_mux[10][17] , \read_value_mux[10][16] , 
        \read_value_mux[10][15] , \read_value_mux[10][14] , 
        \read_value_mux[10][13] , \read_value_mux[10][12] , 
        \read_value_mux[10][11] , \read_value_mux[10][10] , 
        \read_value_mux[10][9] , \read_value_mux[10][8] , 
        \read_value_mux[10][7] , \read_value_mux[10][6] , 
        \read_value_mux[10][5] , \read_value_mux[10][4] , 
        \read_value_mux[10][3] , \read_value_mux[10][2] , 
        \read_value_mux[10][1] , \read_value_mux[10][0] , 
        \read_value_mux[9][31] , \read_value_mux[9][30] , 
        \read_value_mux[9][29] , \read_value_mux[9][28] , 
        \read_value_mux[9][27] , \read_value_mux[9][26] , 
        \read_value_mux[9][25] , \read_value_mux[9][24] , 
        \read_value_mux[9][23] , \read_value_mux[9][22] , 
        \read_value_mux[9][21] , \read_value_mux[9][20] , 
        \read_value_mux[9][19] , \read_value_mux[9][18] , 
        \read_value_mux[9][17] , \read_value_mux[9][16] , 
        \read_value_mux[9][15] , \read_value_mux[9][14] , 
        \read_value_mux[9][13] , \read_value_mux[9][12] , 
        \read_value_mux[9][11] , \read_value_mux[9][10] , 
        \read_value_mux[9][9] , \read_value_mux[9][8] , \read_value_mux[9][7] , 
        \read_value_mux[9][6] , \read_value_mux[9][5] , \read_value_mux[9][4] , 
        \read_value_mux[9][3] , \read_value_mux[9][2] , \read_value_mux[9][1] , 
        \read_value_mux[9][0] , \read_value_mux[8][31] , 
        \read_value_mux[8][30] , \read_value_mux[8][29] , 
        \read_value_mux[8][28] , \read_value_mux[8][27] , 
        \read_value_mux[8][26] , \read_value_mux[8][25] , 
        \read_value_mux[8][24] , \read_value_mux[8][23] , 
        \read_value_mux[8][22] , \read_value_mux[8][21] , 
        \read_value_mux[8][20] , \read_value_mux[8][19] , 
        \read_value_mux[8][18] , \read_value_mux[8][17] , 
        \read_value_mux[8][16] , \read_value_mux[8][15] , 
        \read_value_mux[8][14] , \read_value_mux[8][13] , 
        \read_value_mux[8][12] , \read_value_mux[8][11] , 
        \read_value_mux[8][10] , \read_value_mux[8][9] , 
        \read_value_mux[8][8] , \read_value_mux[8][7] , \read_value_mux[8][6] , 
        \read_value_mux[8][5] , \read_value_mux[8][4] , \read_value_mux[8][3] , 
        \read_value_mux[8][2] , \read_value_mux[8][1] , \read_value_mux[8][0] , 
        \read_value_mux[7][31] , \read_value_mux[7][30] , 
        \read_value_mux[7][29] , \read_value_mux[7][28] , 
        \read_value_mux[7][27] , \read_value_mux[7][26] , 
        \read_value_mux[7][25] , \read_value_mux[7][24] , 
        \read_value_mux[7][23] , \read_value_mux[7][22] , 
        \read_value_mux[7][21] , \read_value_mux[7][20] , 
        \read_value_mux[7][19] , \read_value_mux[7][18] , 
        \read_value_mux[7][17] , \read_value_mux[7][16] , 
        \read_value_mux[7][15] , \read_value_mux[7][14] , 
        \read_value_mux[7][13] , \read_value_mux[7][12] , 
        \read_value_mux[7][11] , \read_value_mux[7][10] , 
        \read_value_mux[7][9] , \read_value_mux[7][8] , \read_value_mux[7][7] , 
        \read_value_mux[7][6] , \read_value_mux[7][5] , \read_value_mux[7][4] , 
        \read_value_mux[7][3] , \read_value_mux[7][2] , \read_value_mux[7][1] , 
        \read_value_mux[7][0] , \read_value_mux[6][31] , 
        \read_value_mux[6][30] , \read_value_mux[6][29] , 
        \read_value_mux[6][28] , \read_value_mux[6][27] , 
        \read_value_mux[6][26] , \read_value_mux[6][25] , 
        \read_value_mux[6][24] , \read_value_mux[6][23] , 
        \read_value_mux[6][22] , \read_value_mux[6][21] , 
        \read_value_mux[6][20] , \read_value_mux[6][19] , 
        \read_value_mux[6][18] , \read_value_mux[6][17] , 
        \read_value_mux[6][16] , \read_value_mux[6][15] , 
        \read_value_mux[6][14] , \read_value_mux[6][13] , 
        \read_value_mux[6][12] , \read_value_mux[6][11] , 
        \read_value_mux[6][10] , \read_value_mux[6][9] , 
        \read_value_mux[6][8] , \read_value_mux[6][7] , \read_value_mux[6][6] , 
        \read_value_mux[6][5] , \read_value_mux[6][4] , \read_value_mux[6][3] , 
        \read_value_mux[6][2] , \read_value_mux[6][1] , \read_value_mux[6][0] , 
        \read_value_mux[5][31] , \read_value_mux[5][30] , 
        \read_value_mux[5][29] , \read_value_mux[5][28] , 
        \read_value_mux[5][27] , \read_value_mux[5][26] , 
        \read_value_mux[5][25] , \read_value_mux[5][24] , 
        \read_value_mux[5][23] , \read_value_mux[5][22] , 
        \read_value_mux[5][21] , \read_value_mux[5][20] , 
        \read_value_mux[5][19] , \read_value_mux[5][18] , 
        \read_value_mux[5][17] , \read_value_mux[5][16] , 
        \read_value_mux[5][15] , \read_value_mux[5][14] , 
        \read_value_mux[5][13] , \read_value_mux[5][12] , 
        \read_value_mux[5][11] , \read_value_mux[5][10] , 
        \read_value_mux[5][9] , \read_value_mux[5][8] , \read_value_mux[5][7] , 
        \read_value_mux[5][6] , \read_value_mux[5][5] , \read_value_mux[5][4] , 
        \read_value_mux[5][3] , \read_value_mux[5][2] , \read_value_mux[5][1] , 
        \read_value_mux[5][0] , \read_value_mux[4][31] , 
        \read_value_mux[4][30] , \read_value_mux[4][29] , 
        \read_value_mux[4][28] , \read_value_mux[4][27] , 
        \read_value_mux[4][26] , \read_value_mux[4][25] , 
        \read_value_mux[4][24] , \read_value_mux[4][23] , 
        \read_value_mux[4][22] , \read_value_mux[4][21] , 
        \read_value_mux[4][20] , \read_value_mux[4][19] , 
        \read_value_mux[4][18] , \read_value_mux[4][17] , 
        \read_value_mux[4][16] , \read_value_mux[4][15] , 
        \read_value_mux[4][14] , \read_value_mux[4][13] , 
        \read_value_mux[4][12] , \read_value_mux[4][11] , 
        \read_value_mux[4][10] , \read_value_mux[4][9] , 
        \read_value_mux[4][8] , \read_value_mux[4][7] , \read_value_mux[4][6] , 
        \read_value_mux[4][5] , \read_value_mux[4][4] , \read_value_mux[4][3] , 
        \read_value_mux[4][2] , \read_value_mux[4][1] , \read_value_mux[4][0] , 
        \read_value_mux[3][31] , \read_value_mux[3][30] , 
        \read_value_mux[3][29] , \read_value_mux[3][28] , 
        \read_value_mux[3][27] , \read_value_mux[3][26] , 
        \read_value_mux[3][25] , \read_value_mux[3][24] , 
        \read_value_mux[3][23] , \read_value_mux[3][22] , 
        \read_value_mux[3][21] , \read_value_mux[3][20] , 
        \read_value_mux[3][19] , \read_value_mux[3][18] , 
        \read_value_mux[3][17] , \read_value_mux[3][16] , 
        \read_value_mux[3][15] , \read_value_mux[3][14] , 
        \read_value_mux[3][13] , \read_value_mux[3][12] , 
        \read_value_mux[3][11] , \read_value_mux[3][10] , 
        \read_value_mux[3][9] , \read_value_mux[3][8] , \read_value_mux[3][7] , 
        \read_value_mux[3][6] , \read_value_mux[3][5] , \read_value_mux[3][4] , 
        \read_value_mux[3][3] , \read_value_mux[3][2] , \read_value_mux[3][1] , 
        \read_value_mux[3][0] , \read_value_mux[2][31] , 
        \read_value_mux[2][30] , \read_value_mux[2][29] , 
        \read_value_mux[2][28] , \read_value_mux[2][27] , 
        \read_value_mux[2][26] , \read_value_mux[2][25] , 
        \read_value_mux[2][24] , \read_value_mux[2][23] , 
        \read_value_mux[2][22] , \read_value_mux[2][21] , 
        \read_value_mux[2][20] , \read_value_mux[2][19] , 
        \read_value_mux[2][18] , \read_value_mux[2][17] , 
        \read_value_mux[2][16] , \read_value_mux[2][15] , 
        \read_value_mux[2][14] , \read_value_mux[2][13] , 
        \read_value_mux[2][12] , \read_value_mux[2][11] , 
        \read_value_mux[2][10] , \read_value_mux[2][9] , 
        \read_value_mux[2][8] , \read_value_mux[2][7] , \read_value_mux[2][6] , 
        \read_value_mux[2][5] , \read_value_mux[2][4] , \read_value_mux[2][3] , 
        \read_value_mux[2][2] , \read_value_mux[2][1] , \read_value_mux[2][0] , 
        \read_value_mux[1][31] , \read_value_mux[1][30] , 
        \read_value_mux[1][29] , \read_value_mux[1][28] , 
        \read_value_mux[1][27] , \read_value_mux[1][26] , 
        \read_value_mux[1][25] , \read_value_mux[1][24] , 
        \read_value_mux[1][23] , \read_value_mux[1][22] , 
        \read_value_mux[1][21] , \read_value_mux[1][20] , 
        \read_value_mux[1][19] , \read_value_mux[1][18] , 
        \read_value_mux[1][17] , \read_value_mux[1][16] , 
        \read_value_mux[1][15] , \read_value_mux[1][14] , 
        \read_value_mux[1][13] , \read_value_mux[1][12] , 
        \read_value_mux[1][11] , \read_value_mux[1][10] , 
        \read_value_mux[1][9] , \read_value_mux[1][8] , \read_value_mux[1][7] , 
        \read_value_mux[1][6] , \read_value_mux[1][5] , \read_value_mux[1][4] , 
        \read_value_mux[1][3] , \read_value_mux[1][2] , \read_value_mux[1][1] , 
        \read_value_mux[1][0] , \read_value_mux[0][31] , 
        \read_value_mux[0][30] , \read_value_mux[0][29] , 
        \read_value_mux[0][28] , \read_value_mux[0][27] , 
        \read_value_mux[0][26] , \read_value_mux[0][25] , 
        \read_value_mux[0][24] , \read_value_mux[0][23] , 
        \read_value_mux[0][22] , \read_value_mux[0][21] , 
        \read_value_mux[0][20] , \read_value_mux[0][19] , 
        \read_value_mux[0][18] , \read_value_mux[0][17] , 
        \read_value_mux[0][16] , \read_value_mux[0][15] , 
        \read_value_mux[0][14] , \read_value_mux[0][13] , 
        \read_value_mux[0][12] , \read_value_mux[0][11] , 
        \read_value_mux[0][10] , \read_value_mux[0][9] , 
        \read_value_mux[0][8] , \read_value_mux[0][7] , \read_value_mux[0][6] , 
        \read_value_mux[0][5] , \read_value_mux[0][4] , \read_value_mux[0][3] , 
        \read_value_mux[0][2] , \read_value_mux[0][1] , \read_value_mux[0][0] }), .select_i(read_index), .data_o(read_value) );
  DFFX1_RVT \words[30]/data_ff/data_reg[31]  ( .D(\words[30]/data_i[31] ), 
        .CLK(clk), .Q(\read_value_mux[30][31] ), .QN(n1674) );
  DFFX1_RVT \words[17]/data_ff/data_reg[31]  ( .D(\words[17]/data_i[31] ), 
        .CLK(clk), .Q(\read_value_mux[17][31] ), .QN(n1673) );
  DFFX1_RVT \words[17]/data_ff/data_reg[0]  ( .D(\words[17]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[17][0] ), .QN(n1672) );
  DFFX1_RVT \words[17]/data_ff/data_reg[29]  ( .D(\words[17]/data_i[29] ), 
        .CLK(clk), .Q(\read_value_mux[17][29] ), .QN(n1671) );
  DFFX1_RVT \words[10]/data_ff/data_reg[31]  ( .D(\words[10]/data_i[31] ), 
        .CLK(clk), .Q(\read_value_mux[10][31] ), .QN(n1670) );
  DFFX1_RVT \words[10]/data_ff/data_reg[29]  ( .D(\words[10]/data_i[29] ), 
        .CLK(clk), .Q(\read_value_mux[10][29] ), .QN(n1669) );
  DFFX1_RVT \words[1]/data_ff/data_reg[31]  ( .D(\words[1]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[1][31] ), .QN(n1668) );
  DFFX1_RVT \words[1]/data_ff/data_reg[0]  ( .D(\words[1]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[1][0] ), .QN(n1667) );
  DFFX1_RVT \words[1]/data_ff/data_reg[29]  ( .D(\words[1]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[1][29] ), .QN(n1666) );
  DFFX1_RVT \words[6]/data_ff/data_reg[31]  ( .D(\words[6]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[6][31] ), .QN(n1665) );
  DFFX1_RVT \words[6]/data_ff/data_reg[0]  ( .D(\words[6]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[6][0] ), .QN(n1664) );
  DFFX1_RVT \words[6]/data_ff/data_reg[29]  ( .D(\words[6]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[6][29] ), .QN(n1663) );
  DFFX1_RVT \words[5]/data_ff/data_reg[31]  ( .D(\words[5]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[5][31] ), .QN(n1662) );
  DFFX1_RVT \words[5]/data_ff/data_reg[29]  ( .D(\words[5]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[5][29] ), .QN(n1661) );
  DFFX1_RVT \words[2]/data_ff/data_reg[31]  ( .D(\words[2]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[2][31] ), .QN(n1660) );
  DFFX1_RVT \words[2]/data_ff/data_reg[0]  ( .D(\words[2]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[2][0] ), .QN(n1659) );
  DFFX1_RVT \words[2]/data_ff/data_reg[29]  ( .D(\words[2]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[2][29] ), .QN(n1658) );
  DFFX1_RVT \words[28]/data_ff/data_reg[31]  ( .D(\words[28]/data_i[31] ), 
        .CLK(clk), .Q(\read_value_mux[28][31] ), .QN(n1657) );
  DFFX1_RVT \words[28]/data_ff/data_reg[29]  ( .D(\words[28]/data_i[29] ), 
        .CLK(clk), .Q(\read_value_mux[28][29] ), .QN(n1656) );
  DFFX1_RVT \words[19]/data_ff/data_reg[31]  ( .D(\words[19]/data_i[31] ), 
        .CLK(clk), .Q(\read_value_mux[19][31] ), .QN(n1655) );
  DFFX1_RVT \words[19]/data_ff/data_reg[29]  ( .D(\words[19]/data_i[29] ), 
        .CLK(clk), .Q(\read_value_mux[19][29] ), .QN(n1654) );
  DFFX1_RVT \words[4]/data_ff/data_reg[31]  ( .D(\words[4]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[4][31] ), .QN(n1653) );
  DFFX1_RVT \words[4]/data_ff/data_reg[0]  ( .D(\words[4]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[4][0] ), .QN(n1652) );
  DFFX1_RVT \words[4]/data_ff/data_reg[29]  ( .D(\words[4]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[4][29] ), .QN(n1651) );
  DFFX1_RVT \words[7]/data_ff/data_reg[31]  ( .D(\words[7]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[7][31] ), .QN(n1650) );
  DFFX1_RVT \words[7]/data_ff/data_reg[29]  ( .D(\words[7]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[7][29] ), .QN(n1649) );
  DFFX1_RVT \words[3]/data_ff/data_reg[31]  ( .D(\words[3]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[3][31] ), .QN(n1648) );
  DFFX1_RVT \words[3]/data_ff/data_reg[0]  ( .D(\words[3]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[3][0] ), .QN(n1647) );
  DFFX1_RVT \words[3]/data_ff/data_reg[29]  ( .D(\words[3]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[3][29] ), .QN(n1646) );
  DFFX1_RVT \words[0]/data_ff/data_reg[31]  ( .D(\words[0]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[0][31] ), .QN(n1645) );
  DFFX1_RVT \words[0]/data_ff/data_reg[0]  ( .D(\words[0]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[0][0] ), .QN(n1644) );
  DFFX1_RVT \words[0]/data_ff/data_reg[29]  ( .D(\words[0]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[0][29] ), .QN(n1643) );
  DFFX1_RVT \words[17]/data_ff/data_reg[28]  ( .D(\words[17]/data_i[28] ), 
        .CLK(clk), .Q(\read_value_mux[17][28] ), .QN(n1642) );
  DFFX1_RVT \words[1]/data_ff/data_reg[28]  ( .D(\words[1]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[1][28] ), .QN(n1641) );
  DFFX1_RVT \words[6]/data_ff/data_reg[28]  ( .D(\words[6]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[6][28] ), .QN(n1640) );
  DFFX1_RVT \words[2]/data_ff/data_reg[28]  ( .D(\words[2]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[2][28] ), .QN(n1639) );
  DFFX1_RVT \words[4]/data_ff/data_reg[28]  ( .D(\words[4]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[4][28] ), .QN(n1638) );
  DFFX1_RVT \words[3]/data_ff/data_reg[28]  ( .D(\words[3]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[3][28] ), .QN(n1637) );
  DFFX1_RVT \words[0]/data_ff/data_reg[28]  ( .D(\words[0]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[0][28] ), .QN(n1636) );
  DFFX1_RVT \words[25]/data_ff/data_reg[31]  ( .D(\words[25]/data_i[31] ), 
        .CLK(clk), .Q(\read_value_mux[25][31] ), .QN(n1629) );
  DFFX1_RVT \words[25]/data_ff/data_reg[0]  ( .D(\words[25]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[25][0] ), .QN(n1628) );
  DFFX1_RVT \words[25]/data_ff/data_reg[29]  ( .D(\words[25]/data_i[29] ), 
        .CLK(clk), .Q(\read_value_mux[25][29] ), .QN(n1627) );
  DFFX1_RVT \words[30]/data_ff/data_reg[0]  ( .D(\words[30]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[30][0] ), .QN(n1626) );
  DFFX1_RVT \words[30]/data_ff/data_reg[29]  ( .D(\words[30]/data_i[29] ), 
        .CLK(clk), .Q(\read_value_mux[30][29] ), .QN(n1625) );
  DFFX1_RVT \words[29]/data_ff/data_reg[31]  ( .D(\words[29]/data_i[31] ), 
        .CLK(clk), .Q(\read_value_mux[29][31] ), .QN(n1624) );
  DFFX1_RVT \words[29]/data_ff/data_reg[0]  ( .D(\words[29]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[29][0] ), .QN(n1623) );
  DFFX1_RVT \words[29]/data_ff/data_reg[29]  ( .D(\words[29]/data_i[29] ), 
        .CLK(clk), .Q(\read_value_mux[29][29] ), .QN(n1622) );
  DFFX1_RVT \words[26]/data_ff/data_reg[31]  ( .D(\words[26]/data_i[31] ), 
        .CLK(clk), .Q(\read_value_mux[26][31] ), .QN(n1621) );
  DFFX1_RVT \words[26]/data_ff/data_reg[0]  ( .D(\words[26]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[26][0] ), .QN(n1620) );
  DFFX1_RVT \words[26]/data_ff/data_reg[29]  ( .D(\words[26]/data_i[29] ), 
        .CLK(clk), .Q(\read_value_mux[26][29] ), .QN(n1619) );
  DFFX1_RVT \words[9]/data_ff/data_reg[28]  ( .D(\words[9]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[9][28] ), .QN(n1618) );
  DFFX1_RVT \words[14]/data_ff/data_reg[31]  ( .D(\words[14]/data_i[31] ), 
        .CLK(clk), .Q(\read_value_mux[14][31] ), .QN(n1617) );
  DFFX1_RVT \words[14]/data_ff/data_reg[0]  ( .D(\words[14]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[14][0] ), .QN(n1616) );
  DFFX1_RVT \words[14]/data_ff/data_reg[29]  ( .D(\words[14]/data_i[29] ), 
        .CLK(clk), .Q(\read_value_mux[14][29] ), .QN(n1615) );
  DFFX1_RVT \words[22]/data_ff/data_reg[31]  ( .D(\words[22]/data_i[31] ), 
        .CLK(clk), .Q(\read_value_mux[22][31] ), .QN(n1614) );
  DFFX1_RVT \words[22]/data_ff/data_reg[0]  ( .D(\words[22]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[22][0] ), .QN(n1613) );
  DFFX1_RVT \words[22]/data_ff/data_reg[29]  ( .D(\words[22]/data_i[29] ), 
        .CLK(clk), .Q(\read_value_mux[22][29] ), .QN(n1612) );
  DFFX1_RVT \words[21]/data_ff/data_reg[31]  ( .D(\words[21]/data_i[31] ), 
        .CLK(clk), .Q(\read_value_mux[21][31] ), .QN(n1611) );
  DFFX1_RVT \words[21]/data_ff/data_reg[0]  ( .D(\words[21]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[21][0] ), .QN(n1610) );
  DFFX1_RVT \words[21]/data_ff/data_reg[29]  ( .D(\words[21]/data_i[29] ), 
        .CLK(clk), .Q(\read_value_mux[21][29] ), .QN(n1609) );
  DFFX1_RVT \words[18]/data_ff/data_reg[31]  ( .D(\words[18]/data_i[31] ), 
        .CLK(clk), .Q(\read_value_mux[18][31] ), .QN(n1608) );
  DFFX1_RVT \words[18]/data_ff/data_reg[0]  ( .D(\words[18]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[18][0] ), .QN(n1607) );
  DFFX1_RVT \words[18]/data_ff/data_reg[29]  ( .D(\words[18]/data_i[29] ), 
        .CLK(clk), .Q(\read_value_mux[18][29] ), .QN(n1606) );
  DFFX1_RVT \words[13]/data_ff/data_reg[31]  ( .D(\words[13]/data_i[31] ), 
        .CLK(clk), .Q(\read_value_mux[13][31] ), .QN(n1605) );
  DFFX1_RVT \words[13]/data_ff/data_reg[0]  ( .D(\words[13]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[13][0] ), .QN(n1604) );
  DFFX1_RVT \words[13]/data_ff/data_reg[29]  ( .D(\words[13]/data_i[29] ), 
        .CLK(clk), .Q(\read_value_mux[13][29] ), .QN(n1603) );
  DFFX1_RVT \words[10]/data_ff/data_reg[0]  ( .D(\words[10]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[10][0] ), .QN(n1602) );
  DFFX1_RVT \words[5]/data_ff/data_reg[0]  ( .D(\words[5]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[5][0] ), .QN(n1601) );
  DFFX1_RVT \words[8]/data_ff/data_reg[31]  ( .D(\words[8]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[8][31] ), .QN(n1600) );
  DFFX1_RVT \words[8]/data_ff/data_reg[0]  ( .D(\words[8]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[8][0] ), .QN(n1599) );
  DFFX1_RVT \words[8]/data_ff/data_reg[29]  ( .D(\words[8]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[8][29] ), .QN(n1598) );
  DFFX1_RVT \words[28]/data_ff/data_reg[0]  ( .D(\words[28]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[28][0] ), .QN(n1597) );
  DFFX1_RVT \words[31]/data_ff/data_reg[31]  ( .D(\words[31]/data_i[31] ), 
        .CLK(clk), .Q(\read_value_mux[31][31] ), .QN(n1596) );
  DFFX1_RVT \words[31]/data_ff/data_reg[0]  ( .D(\words[31]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[31][0] ), .QN(n1595) );
  DFFX1_RVT \words[31]/data_ff/data_reg[29]  ( .D(\words[31]/data_i[29] ), 
        .CLK(clk), .Q(\read_value_mux[31][29] ), .QN(n1594) );
  DFFX1_RVT \words[27]/data_ff/data_reg[31]  ( .D(\words[27]/data_i[31] ), 
        .CLK(clk), .Q(\read_value_mux[27][31] ), .QN(n1593) );
  DFFX1_RVT \words[27]/data_ff/data_reg[0]  ( .D(\words[27]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[27][0] ), .QN(n1592) );
  DFFX1_RVT \words[27]/data_ff/data_reg[29]  ( .D(\words[27]/data_i[29] ), 
        .CLK(clk), .Q(\read_value_mux[27][29] ), .QN(n1591) );
  DFFX1_RVT \words[24]/data_ff/data_reg[31]  ( .D(\words[24]/data_i[31] ), 
        .CLK(clk), .Q(\read_value_mux[24][31] ), .QN(n1590) );
  DFFX1_RVT \words[24]/data_ff/data_reg[0]  ( .D(\words[24]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[24][0] ), .QN(n1589) );
  DFFX1_RVT \words[24]/data_ff/data_reg[29]  ( .D(\words[24]/data_i[29] ), 
        .CLK(clk), .Q(\read_value_mux[24][29] ), .QN(n1588) );
  DFFX1_RVT \words[11]/data_ff/data_reg[31]  ( .D(\words[11]/data_i[31] ), 
        .CLK(clk), .Q(\read_value_mux[11][31] ), .QN(n1587) );
  DFFX1_RVT \words[11]/data_ff/data_reg[0]  ( .D(\words[11]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[11][0] ), .QN(n1586) );
  DFFX1_RVT \words[11]/data_ff/data_reg[29]  ( .D(\words[11]/data_i[29] ), 
        .CLK(clk), .Q(\read_value_mux[11][29] ), .QN(n1585) );
  DFFX1_RVT \words[15]/data_ff/data_reg[31]  ( .D(\words[15]/data_i[31] ), 
        .CLK(clk), .Q(\read_value_mux[15][31] ), .QN(n1584) );
  DFFX1_RVT \words[15]/data_ff/data_reg[0]  ( .D(\words[15]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[15][0] ), .QN(n1583) );
  DFFX1_RVT \words[15]/data_ff/data_reg[29]  ( .D(\words[15]/data_i[29] ), 
        .CLK(clk), .Q(\read_value_mux[15][29] ), .QN(n1582) );
  DFFX1_RVT \words[20]/data_ff/data_reg[31]  ( .D(\words[20]/data_i[31] ), 
        .CLK(clk), .Q(\read_value_mux[20][31] ), .QN(n1581) );
  DFFX1_RVT \words[20]/data_ff/data_reg[0]  ( .D(\words[20]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[20][0] ), .QN(n1580) );
  DFFX1_RVT \words[20]/data_ff/data_reg[29]  ( .D(\words[20]/data_i[29] ), 
        .CLK(clk), .Q(\read_value_mux[20][29] ), .QN(n1579) );
  DFFX1_RVT \words[23]/data_ff/data_reg[31]  ( .D(\words[23]/data_i[31] ), 
        .CLK(clk), .Q(\read_value_mux[23][31] ), .QN(n1578) );
  DFFX1_RVT \words[23]/data_ff/data_reg[0]  ( .D(\words[23]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[23][0] ), .QN(n1577) );
  DFFX1_RVT \words[23]/data_ff/data_reg[29]  ( .D(\words[23]/data_i[29] ), 
        .CLK(clk), .Q(\read_value_mux[23][29] ), .QN(n1576) );
  DFFX1_RVT \words[19]/data_ff/data_reg[0]  ( .D(\words[19]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[19][0] ), .QN(n1575) );
  DFFX1_RVT \words[16]/data_ff/data_reg[31]  ( .D(\words[16]/data_i[31] ), 
        .CLK(clk), .Q(\read_value_mux[16][31] ), .QN(n1574) );
  DFFX1_RVT \words[16]/data_ff/data_reg[0]  ( .D(\words[16]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[16][0] ), .QN(n1573) );
  DFFX1_RVT \words[16]/data_ff/data_reg[29]  ( .D(\words[16]/data_i[29] ), 
        .CLK(clk), .Q(\read_value_mux[16][29] ), .QN(n1572) );
  DFFX1_RVT \words[12]/data_ff/data_reg[31]  ( .D(\words[12]/data_i[31] ), 
        .CLK(clk), .Q(\read_value_mux[12][31] ), .QN(n1571) );
  DFFX1_RVT \words[12]/data_ff/data_reg[0]  ( .D(\words[12]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[12][0] ), .QN(n1570) );
  DFFX1_RVT \words[12]/data_ff/data_reg[29]  ( .D(\words[12]/data_i[29] ), 
        .CLK(clk), .Q(\read_value_mux[12][29] ), .QN(n1569) );
  DFFX1_RVT \words[7]/data_ff/data_reg[0]  ( .D(\words[7]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[7][0] ), .QN(n1568) );
  DFFX1_RVT \words[25]/data_ff/data_reg[28]  ( .D(\words[25]/data_i[28] ), 
        .CLK(clk), .Q(\read_value_mux[25][28] ), .QN(n1567) );
  DFFX1_RVT \words[30]/data_ff/data_reg[28]  ( .D(\words[30]/data_i[28] ), 
        .CLK(clk), .Q(\read_value_mux[30][28] ), .QN(n1566) );
  DFFX1_RVT \words[29]/data_ff/data_reg[28]  ( .D(\words[29]/data_i[28] ), 
        .CLK(clk), .Q(\read_value_mux[29][28] ), .QN(n1565) );
  DFFX1_RVT \words[26]/data_ff/data_reg[28]  ( .D(\words[26]/data_i[28] ), 
        .CLK(clk), .Q(\read_value_mux[26][28] ), .QN(n1564) );
  DFFX1_RVT \words[14]/data_ff/data_reg[28]  ( .D(\words[14]/data_i[28] ), 
        .CLK(clk), .Q(\read_value_mux[14][28] ), .QN(n1563) );
  DFFX1_RVT \words[22]/data_ff/data_reg[28]  ( .D(\words[22]/data_i[28] ), 
        .CLK(clk), .Q(\read_value_mux[22][28] ), .QN(n1562) );
  DFFX1_RVT \words[21]/data_ff/data_reg[28]  ( .D(\words[21]/data_i[28] ), 
        .CLK(clk), .Q(\read_value_mux[21][28] ), .QN(n1561) );
  DFFX1_RVT \words[18]/data_ff/data_reg[28]  ( .D(\words[18]/data_i[28] ), 
        .CLK(clk), .Q(\read_value_mux[18][28] ), .QN(n1560) );
  DFFX1_RVT \words[13]/data_ff/data_reg[28]  ( .D(\words[13]/data_i[28] ), 
        .CLK(clk), .Q(\read_value_mux[13][28] ), .QN(n1559) );
  DFFX1_RVT \words[10]/data_ff/data_reg[28]  ( .D(\words[10]/data_i[28] ), 
        .CLK(clk), .Q(\read_value_mux[10][28] ), .QN(n1558) );
  DFFX1_RVT \words[5]/data_ff/data_reg[28]  ( .D(\words[5]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[5][28] ), .QN(n1557) );
  DFFX1_RVT \words[8]/data_ff/data_reg[28]  ( .D(\words[8]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[8][28] ), .QN(n1556) );
  DFFX1_RVT \words[28]/data_ff/data_reg[28]  ( .D(\words[28]/data_i[28] ), 
        .CLK(clk), .Q(\read_value_mux[28][28] ), .QN(n1555) );
  DFFX1_RVT \words[31]/data_ff/data_reg[28]  ( .D(\words[31]/data_i[28] ), 
        .CLK(clk), .Q(\read_value_mux[31][28] ), .QN(n1554) );
  DFFX1_RVT \words[27]/data_ff/data_reg[28]  ( .D(\words[27]/data_i[28] ), 
        .CLK(clk), .Q(\read_value_mux[27][28] ), .QN(n1553) );
  DFFX1_RVT \words[24]/data_ff/data_reg[28]  ( .D(\words[24]/data_i[28] ), 
        .CLK(clk), .Q(\read_value_mux[24][28] ), .QN(n1552) );
  DFFX1_RVT \words[11]/data_ff/data_reg[28]  ( .D(\words[11]/data_i[28] ), 
        .CLK(clk), .Q(\read_value_mux[11][28] ), .QN(n1551) );
  DFFX1_RVT \words[15]/data_ff/data_reg[28]  ( .D(\words[15]/data_i[28] ), 
        .CLK(clk), .Q(\read_value_mux[15][28] ), .QN(n1550) );
  DFFX1_RVT \words[20]/data_ff/data_reg[28]  ( .D(\words[20]/data_i[28] ), 
        .CLK(clk), .Q(\read_value_mux[20][28] ), .QN(n1549) );
  DFFX1_RVT \words[23]/data_ff/data_reg[28]  ( .D(\words[23]/data_i[28] ), 
        .CLK(clk), .Q(\read_value_mux[23][28] ), .QN(n1548) );
  DFFX1_RVT \words[19]/data_ff/data_reg[28]  ( .D(\words[19]/data_i[28] ), 
        .CLK(clk), .Q(\read_value_mux[19][28] ), .QN(n1547) );
  DFFX1_RVT \words[16]/data_ff/data_reg[28]  ( .D(\words[16]/data_i[28] ), 
        .CLK(clk), .Q(\read_value_mux[16][28] ), .QN(n1546) );
  DFFX1_RVT \words[12]/data_ff/data_reg[28]  ( .D(\words[12]/data_i[28] ), 
        .CLK(clk), .Q(\read_value_mux[12][28] ), .QN(n1545) );
  DFFX1_RVT \words[7]/data_ff/data_reg[28]  ( .D(\words[7]/data_i[28] ), .CLK(
        clk), .Q(\read_value_mux[7][28] ), .QN(n1544) );
  DFFX1_RVT \words[7]/data_ff/data_reg[1]  ( .D(\words[7]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[7][1] ), .QN(n28) );
  DFFX1_RVT \words[6]/data_ff/data_reg[1]  ( .D(\words[6]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[6][1] ), .QN(n26) );
  DFFX1_RVT \words[5]/data_ff/data_reg[1]  ( .D(\words[5]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[5][1] ), .QN(n23) );
  DFFX1_RVT \words[4]/data_ff/data_reg[1]  ( .D(\words[4]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[4][1] ), .QN(n21) );
  DFFX1_RVT \words[3]/data_ff/data_reg[1]  ( .D(\words[3]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[3][1] ), .QN(n18) );
  DFFX1_RVT \words[30]/data_ff/data_reg[1]  ( .D(\words[30]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[30][1] ), .QN(n88) );
  DFFX1_RVT \words[2]/data_ff/data_reg[1]  ( .D(\words[2]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[2][1] ), .QN(n16) );
  DFFX1_RVT \words[28]/data_ff/data_reg[1]  ( .D(\words[28]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[28][1] ), .QN(n83) );
  DFFX1_RVT \words[23]/data_ff/data_reg[1]  ( .D(\words[23]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[23][1] ), .QN(n71) );
  DFFX1_RVT \words[1]/data_ff/data_reg[1]  ( .D(\words[1]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[1][1] ), .QN(n14) );
  DFFX1_RVT \words[19]/data_ff/data_reg[1]  ( .D(\words[19]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[19][1] ), .QN(n60) );
  DFFX1_RVT \words[17]/data_ff/data_reg[1]  ( .D(\words[17]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[17][1] ), .QN(n55) );
  DFFX1_RVT \words[12]/data_ff/data_reg[1]  ( .D(\words[12]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[12][1] ), .QN(n43) );
  DFFX1_RVT \words[10]/data_ff/data_reg[1]  ( .D(\words[10]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[10][1] ), .QN(n37) );
  DFFX1_RVT \words[0]/data_ff/data_reg[1]  ( .D(\words[0]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[0][1] ), .QN(n11) );
  DFFX1_RVT \words[6]/data_ff/data_reg[30]  ( .D(\words[6]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[6][30] ), .QN(n27) );
  DFFX1_RVT \words[4]/data_ff/data_reg[30]  ( .D(\words[4]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[4][30] ), .QN(n22) );
  DFFX1_RVT \words[3]/data_ff/data_reg[30]  ( .D(\words[3]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[3][30] ), .QN(n19) );
  DFFX1_RVT \words[2]/data_ff/data_reg[30]  ( .D(\words[2]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[2][30] ), .QN(n17) );
  DFFX1_RVT \words[1]/data_ff/data_reg[30]  ( .D(\words[1]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[1][30] ), .QN(n15) );
  DFFX1_RVT \words[19]/data_ff/data_reg[30]  ( .D(\words[19]/data_i[30] ), 
        .CLK(clk), .Q(\read_value_mux[19][30] ), .QN(n61) );
  DFFX1_RVT \words[17]/data_ff/data_reg[30]  ( .D(\words[17]/data_i[30] ), 
        .CLK(clk), .Q(\read_value_mux[17][30] ), .QN(n56) );
  DFFX1_RVT \words[0]/data_ff/data_reg[30]  ( .D(\words[0]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[0][30] ), .QN(n12) );
  DFFX1_RVT \words[9]/data_ff/data_reg[30]  ( .D(\words[9]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[9][30] ), .QN(n34) );
  DFFX1_RVT \words[8]/data_ff/data_reg[1]  ( .D(\words[8]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[8][1] ), .QN(n30) );
  DFFX1_RVT \words[31]/data_ff/data_reg[1]  ( .D(\words[31]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[31][1] ), .QN(n6) );
  DFFX1_RVT \words[29]/data_ff/data_reg[1]  ( .D(\words[29]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[29][1] ), .QN(n85) );
  DFFX1_RVT \words[27]/data_ff/data_reg[1]  ( .D(\words[27]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[27][1] ), .QN(n81) );
  DFFX1_RVT \words[26]/data_ff/data_reg[1]  ( .D(\words[26]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[26][1] ), .QN(n79) );
  DFFX1_RVT \words[25]/data_ff/data_reg[1]  ( .D(\words[25]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[25][1] ), .QN(n76) );
  DFFX1_RVT \words[24]/data_ff/data_reg[1]  ( .D(\words[24]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[24][1] ), .QN(n74) );
  DFFX1_RVT \words[22]/data_ff/data_reg[1]  ( .D(\words[22]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[22][1] ), .QN(n69) );
  DFFX1_RVT \words[21]/data_ff/data_reg[1]  ( .D(\words[21]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[21][1] ), .QN(n66) );
  DFFX1_RVT \words[20]/data_ff/data_reg[1]  ( .D(\words[20]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[20][1] ), .QN(n64) );
  DFFX1_RVT \words[18]/data_ff/data_reg[1]  ( .D(\words[18]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[18][1] ), .QN(n58) );
  DFFX1_RVT \words[16]/data_ff/data_reg[1]  ( .D(\words[16]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[16][1] ), .QN(n53) );
  DFFX1_RVT \words[15]/data_ff/data_reg[1]  ( .D(\words[15]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[15][1] ), .QN(n50) );
  DFFX1_RVT \words[14]/data_ff/data_reg[1]  ( .D(\words[14]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[14][1] ), .QN(n48) );
  DFFX1_RVT \words[13]/data_ff/data_reg[1]  ( .D(\words[13]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[13][1] ), .QN(n45) );
  DFFX1_RVT \words[11]/data_ff/data_reg[1]  ( .D(\words[11]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[11][1] ), .QN(n39) );
  DFFX1_RVT \words[8]/data_ff/data_reg[30]  ( .D(\words[8]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[8][30] ), .QN(n31) );
  DFFX1_RVT \words[7]/data_ff/data_reg[30]  ( .D(\words[7]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[7][30] ), .QN(n29) );
  DFFX1_RVT \words[5]/data_ff/data_reg[30]  ( .D(\words[5]/data_i[30] ), .CLK(
        clk), .Q(\read_value_mux[5][30] ), .QN(n24) );
  DFFX1_RVT \words[31]/data_ff/data_reg[30]  ( .D(\words[31]/data_i[30] ), 
        .CLK(clk), .Q(\read_value_mux[31][30] ), .QN(n7) );
  DFFX1_RVT \words[30]/data_ff/data_reg[30]  ( .D(\words[30]/data_i[30] ), 
        .CLK(clk), .Q(\read_value_mux[30][30] ), .QN(n89) );
  DFFX1_RVT \words[29]/data_ff/data_reg[30]  ( .D(\words[29]/data_i[30] ), 
        .CLK(clk), .Q(\read_value_mux[29][30] ), .QN(n86) );
  DFFX1_RVT \words[28]/data_ff/data_reg[30]  ( .D(\words[28]/data_i[30] ), 
        .CLK(clk), .Q(\read_value_mux[28][30] ), .QN(n84) );
  DFFX1_RVT \words[27]/data_ff/data_reg[30]  ( .D(\words[27]/data_i[30] ), 
        .CLK(clk), .Q(\read_value_mux[27][30] ), .QN(n82) );
  DFFX1_RVT \words[26]/data_ff/data_reg[30]  ( .D(\words[26]/data_i[30] ), 
        .CLK(clk), .Q(\read_value_mux[26][30] ), .QN(n80) );
  DFFX1_RVT \words[25]/data_ff/data_reg[30]  ( .D(\words[25]/data_i[30] ), 
        .CLK(clk), .Q(\read_value_mux[25][30] ), .QN(n77) );
  DFFX1_RVT \words[24]/data_ff/data_reg[30]  ( .D(\words[24]/data_i[30] ), 
        .CLK(clk), .Q(\read_value_mux[24][30] ), .QN(n75) );
  DFFX1_RVT \words[23]/data_ff/data_reg[30]  ( .D(\words[23]/data_i[30] ), 
        .CLK(clk), .Q(\read_value_mux[23][30] ), .QN(n72) );
  DFFX1_RVT \words[22]/data_ff/data_reg[30]  ( .D(\words[22]/data_i[30] ), 
        .CLK(clk), .Q(\read_value_mux[22][30] ), .QN(n70) );
  DFFX1_RVT \words[21]/data_ff/data_reg[30]  ( .D(\words[21]/data_i[30] ), 
        .CLK(clk), .Q(\read_value_mux[21][30] ), .QN(n67) );
  DFFX1_RVT \words[20]/data_ff/data_reg[30]  ( .D(\words[20]/data_i[30] ), 
        .CLK(clk), .Q(\read_value_mux[20][30] ), .QN(n65) );
  DFFX1_RVT \words[18]/data_ff/data_reg[30]  ( .D(\words[18]/data_i[30] ), 
        .CLK(clk), .Q(\read_value_mux[18][30] ), .QN(n59) );
  DFFX1_RVT \words[16]/data_ff/data_reg[30]  ( .D(\words[16]/data_i[30] ), 
        .CLK(clk), .Q(\read_value_mux[16][30] ), .QN(n54) );
  DFFX1_RVT \words[15]/data_ff/data_reg[30]  ( .D(\words[15]/data_i[30] ), 
        .CLK(clk), .Q(\read_value_mux[15][30] ), .QN(n51) );
  DFFX1_RVT \words[14]/data_ff/data_reg[30]  ( .D(\words[14]/data_i[30] ), 
        .CLK(clk), .Q(\read_value_mux[14][30] ), .QN(n49) );
  DFFX1_RVT \words[13]/data_ff/data_reg[30]  ( .D(\words[13]/data_i[30] ), 
        .CLK(clk), .Q(\read_value_mux[13][30] ), .QN(n46) );
  DFFX1_RVT \words[12]/data_ff/data_reg[30]  ( .D(\words[12]/data_i[30] ), 
        .CLK(clk), .Q(\read_value_mux[12][30] ), .QN(n44) );
  DFFX1_RVT \words[11]/data_ff/data_reg[30]  ( .D(\words[11]/data_i[30] ), 
        .CLK(clk), .Q(\read_value_mux[11][30] ), .QN(n40) );
  DFFX1_RVT \words[10]/data_ff/data_reg[30]  ( .D(\words[10]/data_i[30] ), 
        .CLK(clk), .Q(\read_value_mux[10][30] ), .QN(n38) );
  DFFX1_RVT \words[4]/valid_ff/data_reg[0]  ( .D(\words[4]/valid_i ), .CLK(clk), .Q(\words[4]/valid_o ) );
  DFFX1_RVT \words[6]/valid_ff/data_reg[0]  ( .D(\words[6]/valid_i ), .CLK(clk), .Q(\words[6]/valid_o ) );
  DFFX1_RVT \words[12]/valid_ff/data_reg[0]  ( .D(\words[12]/valid_i ), .CLK(
        clk), .Q(\words[12]/valid_o ) );
  DFFX1_RVT \words[14]/valid_ff/data_reg[0]  ( .D(\words[14]/valid_i ), .CLK(
        clk), .Q(\words[14]/valid_o ) );
  DFFX1_RVT \words[2]/valid_ff/data_reg[0]  ( .D(\words[2]/valid_i ), .CLK(clk), .Q(\words[2]/valid_o ) );
  DFFX1_RVT \words[10]/valid_ff/data_reg[0]  ( .D(\words[10]/valid_i ), .CLK(
        clk), .Q(\words[10]/valid_o ) );
  DFFX1_RVT \words[31]/valid_ff/data_reg[0]  ( .D(\words[31]/valid_i ), .CLK(
        clk), .Q(\words[31]/valid_o ) );
  DFFX1_RVT \words[16]/valid_ff/data_reg[0]  ( .D(\words[16]/valid_i ), .CLK(
        clk), .Q(\words[16]/valid_o ) );
  DFFX1_RVT \words[17]/valid_ff/data_reg[0]  ( .D(\words[17]/valid_i ), .CLK(
        clk), .Q(\words[17]/valid_o ) );
  DFFX1_RVT \words[20]/valid_ff/data_reg[0]  ( .D(\words[20]/valid_i ), .CLK(
        clk), .Q(\words[20]/valid_o ) );
  DFFX1_RVT \words[21]/valid_ff/data_reg[0]  ( .D(\words[21]/valid_i ), .CLK(
        clk), .Q(\words[21]/valid_o ) );
  DFFX1_RVT \words[24]/valid_ff/data_reg[0]  ( .D(\words[24]/valid_i ), .CLK(
        clk), .Q(\words[24]/valid_o ) );
  DFFX1_RVT \words[25]/valid_ff/data_reg[0]  ( .D(\words[25]/valid_i ), .CLK(
        clk), .Q(\words[25]/valid_o ) );
  DFFX1_RVT \words[30]/valid_ff/data_reg[0]  ( .D(\words[30]/valid_i ), .CLK(
        clk), .Q(\words[30]/valid_o ) );
  DFFX1_RVT \words[0]/valid_ff/data_reg[0]  ( .D(\words[0]/valid_i ), .CLK(clk), .Q(\words[0]/valid_o ) );
  DFFX1_RVT \words[8]/valid_ff/data_reg[0]  ( .D(\words[8]/valid_i ), .CLK(clk), .Q(\words[8]/valid_o ) );
  DFFX1_RVT \words[1]/valid_ff/data_reg[0]  ( .D(\words[1]/valid_i ), .CLK(clk), .Q(\words[1]/valid_o ) );
  DFFX1_RVT \words[9]/valid_ff/data_reg[0]  ( .D(\words[9]/valid_i ), .CLK(clk), .Q(\words[9]/valid_o ) );
  DFFX1_RVT \words[5]/valid_ff/data_reg[0]  ( .D(\words[5]/valid_i ), .CLK(clk), .Q(\words[5]/valid_o ) );
  DFFX1_RVT \words[13]/valid_ff/data_reg[0]  ( .D(\words[13]/valid_i ), .CLK(
        clk), .Q(\words[13]/valid_o ) );
  DFFX1_RVT \words[7]/valid_ff/data_reg[0]  ( .D(\words[7]/valid_i ), .CLK(clk), .Q(\words[7]/valid_o ) );
  DFFX1_RVT \words[15]/valid_ff/data_reg[0]  ( .D(\words[15]/valid_i ), .CLK(
        clk), .Q(\words[15]/valid_o ) );
  DFFX1_RVT \words[3]/valid_ff/data_reg[0]  ( .D(\words[3]/valid_i ), .CLK(clk), .Q(\words[3]/valid_o ) );
  DFFX1_RVT \words[11]/valid_ff/data_reg[0]  ( .D(\words[11]/valid_i ), .CLK(
        clk), .Q(\words[11]/valid_o ) );
  DFFX1_RVT \words[18]/valid_ff/data_reg[0]  ( .D(\words[18]/valid_i ), .CLK(
        clk), .Q(\words[18]/valid_o ) );
  DFFX1_RVT \words[19]/valid_ff/data_reg[0]  ( .D(\words[19]/valid_i ), .CLK(
        clk), .Q(\words[19]/valid_o ) );
  DFFX1_RVT \words[22]/valid_ff/data_reg[0]  ( .D(\words[22]/valid_i ), .CLK(
        clk), .Q(\words[22]/valid_o ) );
  DFFX1_RVT \words[23]/valid_ff/data_reg[0]  ( .D(\words[23]/valid_i ), .CLK(
        clk), .Q(\words[23]/valid_o ) );
  DFFX1_RVT \words[26]/valid_ff/data_reg[0]  ( .D(\words[26]/valid_i ), .CLK(
        clk), .Q(\words[26]/valid_o ) );
  DFFX1_RVT \words[27]/valid_ff/data_reg[0]  ( .D(\words[27]/valid_i ), .CLK(
        clk), .Q(\words[27]/valid_o ) );
  DFFX1_RVT \words[28]/valid_ff/data_reg[0]  ( .D(\words[28]/valid_i ), .CLK(
        clk), .Q(\words[28]/valid_o ) );
  DFFX1_RVT \words[29]/valid_ff/data_reg[0]  ( .D(\words[29]/valid_i ), .CLK(
        clk), .Q(\words[29]/valid_o ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[2]  ( .D(\words[1]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[1][2] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[4]  ( .D(\words[1]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[1][4] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[6]  ( .D(\words[1]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[1][6] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[8]  ( .D(\words[1]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[1][8] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[10]  ( .D(\words[1]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[1][10] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[12]  ( .D(\words[1]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[1][12] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[14]  ( .D(\words[1]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[1][14] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[16]  ( .D(\words[1]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[1][16] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[18]  ( .D(\words[1]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[1][18] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[20]  ( .D(\words[1]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[1][20] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[22]  ( .D(\words[1]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[1][22] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[24]  ( .D(\words[1]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[1][24] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[26]  ( .D(\words[1]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[1][26] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[2]  ( .D(\words[2]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[2][2] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[4]  ( .D(\words[2]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[2][4] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[6]  ( .D(\words[2]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[2][6] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[8]  ( .D(\words[2]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[2][8] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[10]  ( .D(\words[2]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[2][10] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[12]  ( .D(\words[2]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[2][12] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[14]  ( .D(\words[2]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[2][14] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[16]  ( .D(\words[2]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[2][16] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[18]  ( .D(\words[2]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[2][18] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[20]  ( .D(\words[2]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[2][20] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[22]  ( .D(\words[2]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[2][22] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[24]  ( .D(\words[2]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[2][24] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[26]  ( .D(\words[2]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[2][26] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[2]  ( .D(\words[5]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[5][2] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[6]  ( .D(\words[5]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[5][6] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[10]  ( .D(\words[5]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[5][10] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[18]  ( .D(\words[5]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[5][18] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[2]  ( .D(\words[6]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[6][2] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[4]  ( .D(\words[6]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[6][4] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[6]  ( .D(\words[6]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[6][6] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[8]  ( .D(\words[6]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[6][8] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[10]  ( .D(\words[6]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[6][10] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[12]  ( .D(\words[6]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[6][12] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[14]  ( .D(\words[6]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[6][14] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[16]  ( .D(\words[6]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[6][16] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[18]  ( .D(\words[6]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[6][18] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[20]  ( .D(\words[6]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[6][20] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[22]  ( .D(\words[6]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[6][22] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[24]  ( .D(\words[6]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[6][24] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[26]  ( .D(\words[6]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[6][26] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[2]  ( .D(\words[17]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[17][2] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[4]  ( .D(\words[17]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[17][4] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[6]  ( .D(\words[17]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[17][6] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[8]  ( .D(\words[17]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[17][8] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[10]  ( .D(\words[17]/data_i[10] ), 
        .CLK(clk), .Q(\read_value_mux[17][10] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[12]  ( .D(\words[17]/data_i[12] ), 
        .CLK(clk), .Q(\read_value_mux[17][12] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[14]  ( .D(\words[17]/data_i[14] ), 
        .CLK(clk), .Q(\read_value_mux[17][14] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[16]  ( .D(\words[17]/data_i[16] ), 
        .CLK(clk), .Q(\read_value_mux[17][16] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[18]  ( .D(\words[17]/data_i[18] ), 
        .CLK(clk), .Q(\read_value_mux[17][18] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[20]  ( .D(\words[17]/data_i[20] ), 
        .CLK(clk), .Q(\read_value_mux[17][20] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[22]  ( .D(\words[17]/data_i[22] ), 
        .CLK(clk), .Q(\read_value_mux[17][22] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[24]  ( .D(\words[17]/data_i[24] ), 
        .CLK(clk), .Q(\read_value_mux[17][24] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[26]  ( .D(\words[17]/data_i[26] ), 
        .CLK(clk), .Q(\read_value_mux[17][26] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[3]  ( .D(\words[1]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[1][3] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[5]  ( .D(\words[1]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[1][5] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[7]  ( .D(\words[1]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[1][7] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[9]  ( .D(\words[1]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[1][9] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[11]  ( .D(\words[1]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[1][11] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[13]  ( .D(\words[1]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[1][13] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[15]  ( .D(\words[1]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[1][15] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[17]  ( .D(\words[1]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[1][17] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[19]  ( .D(\words[1]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[1][19] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[21]  ( .D(\words[1]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[1][21] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[23]  ( .D(\words[1]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[1][23] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[25]  ( .D(\words[1]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[1][25] ) );
  DFFX1_RVT \words[1]/data_ff/data_reg[27]  ( .D(\words[1]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[1][27] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[3]  ( .D(\words[2]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[2][3] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[5]  ( .D(\words[2]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[2][5] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[7]  ( .D(\words[2]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[2][7] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[9]  ( .D(\words[2]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[2][9] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[11]  ( .D(\words[2]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[2][11] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[13]  ( .D(\words[2]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[2][13] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[15]  ( .D(\words[2]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[2][15] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[17]  ( .D(\words[2]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[2][17] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[19]  ( .D(\words[2]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[2][19] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[21]  ( .D(\words[2]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[2][21] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[23]  ( .D(\words[2]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[2][23] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[25]  ( .D(\words[2]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[2][25] ) );
  DFFX1_RVT \words[2]/data_ff/data_reg[27]  ( .D(\words[2]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[2][27] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[3]  ( .D(\words[5]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[5][3] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[7]  ( .D(\words[5]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[5][7] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[11]  ( .D(\words[5]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[5][11] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[19]  ( .D(\words[5]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[5][19] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[27]  ( .D(\words[5]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[5][27] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[3]  ( .D(\words[6]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[6][3] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[5]  ( .D(\words[6]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[6][5] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[7]  ( .D(\words[6]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[6][7] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[9]  ( .D(\words[6]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[6][9] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[11]  ( .D(\words[6]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[6][11] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[13]  ( .D(\words[6]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[6][13] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[15]  ( .D(\words[6]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[6][15] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[17]  ( .D(\words[6]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[6][17] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[19]  ( .D(\words[6]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[6][19] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[21]  ( .D(\words[6]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[6][21] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[23]  ( .D(\words[6]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[6][23] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[25]  ( .D(\words[6]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[6][25] ) );
  DFFX1_RVT \words[6]/data_ff/data_reg[27]  ( .D(\words[6]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[6][27] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[5]  ( .D(\words[10]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[10][5] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[13]  ( .D(\words[10]/data_i[13] ), 
        .CLK(clk), .Q(\read_value_mux[10][13] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[3]  ( .D(\words[17]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[17][3] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[5]  ( .D(\words[17]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[17][5] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[7]  ( .D(\words[17]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[17][7] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[9]  ( .D(\words[17]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[17][9] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[11]  ( .D(\words[17]/data_i[11] ), 
        .CLK(clk), .Q(\read_value_mux[17][11] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[13]  ( .D(\words[17]/data_i[13] ), 
        .CLK(clk), .Q(\read_value_mux[17][13] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[15]  ( .D(\words[17]/data_i[15] ), 
        .CLK(clk), .Q(\read_value_mux[17][15] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[17]  ( .D(\words[17]/data_i[17] ), 
        .CLK(clk), .Q(\read_value_mux[17][17] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[19]  ( .D(\words[17]/data_i[19] ), 
        .CLK(clk), .Q(\read_value_mux[17][19] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[21]  ( .D(\words[17]/data_i[21] ), 
        .CLK(clk), .Q(\read_value_mux[17][21] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[23]  ( .D(\words[17]/data_i[23] ), 
        .CLK(clk), .Q(\read_value_mux[17][23] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[25]  ( .D(\words[17]/data_i[25] ), 
        .CLK(clk), .Q(\read_value_mux[17][25] ) );
  DFFX1_RVT \words[17]/data_ff/data_reg[27]  ( .D(\words[17]/data_i[27] ), 
        .CLK(clk), .Q(\read_value_mux[17][27] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[2]  ( .D(\words[0]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[0][2] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[4]  ( .D(\words[0]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[0][4] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[6]  ( .D(\words[0]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[0][6] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[8]  ( .D(\words[0]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[0][8] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[10]  ( .D(\words[0]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[0][10] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[12]  ( .D(\words[0]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[0][12] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[14]  ( .D(\words[0]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[0][14] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[16]  ( .D(\words[0]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[0][16] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[18]  ( .D(\words[0]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[0][18] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[20]  ( .D(\words[0]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[0][20] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[22]  ( .D(\words[0]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[0][22] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[24]  ( .D(\words[0]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[0][24] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[26]  ( .D(\words[0]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[0][26] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[2]  ( .D(\words[3]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[3][2] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[4]  ( .D(\words[3]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[3][4] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[6]  ( .D(\words[3]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[3][6] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[8]  ( .D(\words[3]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[3][8] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[10]  ( .D(\words[3]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[3][10] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[12]  ( .D(\words[3]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[3][12] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[14]  ( .D(\words[3]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[3][14] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[16]  ( .D(\words[3]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[3][16] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[18]  ( .D(\words[3]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[3][18] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[20]  ( .D(\words[3]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[3][20] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[22]  ( .D(\words[3]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[3][22] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[24]  ( .D(\words[3]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[3][24] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[26]  ( .D(\words[3]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[3][26] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[2]  ( .D(\words[4]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[4][2] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[4]  ( .D(\words[4]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[4][4] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[6]  ( .D(\words[4]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[4][6] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[8]  ( .D(\words[4]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[4][8] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[10]  ( .D(\words[4]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[4][10] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[12]  ( .D(\words[4]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[4][12] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[14]  ( .D(\words[4]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[4][14] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[16]  ( .D(\words[4]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[4][16] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[18]  ( .D(\words[4]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[4][18] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[20]  ( .D(\words[4]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[4][20] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[22]  ( .D(\words[4]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[4][22] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[24]  ( .D(\words[4]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[4][24] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[26]  ( .D(\words[4]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[4][26] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[2]  ( .D(\words[7]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[7][2] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[6]  ( .D(\words[7]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[7][6] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[10]  ( .D(\words[7]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[7][10] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[18]  ( .D(\words[7]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[7][18] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[26]  ( .D(\words[7]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[7][26] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[2]  ( .D(\words[19]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[19][2] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[4]  ( .D(\words[19]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[19][4] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[6]  ( .D(\words[19]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[19][6] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[8]  ( .D(\words[19]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[19][8] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[10]  ( .D(\words[19]/data_i[10] ), 
        .CLK(clk), .Q(\read_value_mux[19][10] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[12]  ( .D(\words[19]/data_i[12] ), 
        .CLK(clk), .Q(\read_value_mux[19][12] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[14]  ( .D(\words[19]/data_i[14] ), 
        .CLK(clk), .Q(\read_value_mux[19][14] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[16]  ( .D(\words[19]/data_i[16] ), 
        .CLK(clk), .Q(\read_value_mux[19][16] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[18]  ( .D(\words[19]/data_i[18] ), 
        .CLK(clk), .Q(\read_value_mux[19][18] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[20]  ( .D(\words[19]/data_i[20] ), 
        .CLK(clk), .Q(\read_value_mux[19][20] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[22]  ( .D(\words[19]/data_i[22] ), 
        .CLK(clk), .Q(\read_value_mux[19][22] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[24]  ( .D(\words[19]/data_i[24] ), 
        .CLK(clk), .Q(\read_value_mux[19][24] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[26]  ( .D(\words[19]/data_i[26] ), 
        .CLK(clk), .Q(\read_value_mux[19][26] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[2]  ( .D(\words[28]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[28][2] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[4]  ( .D(\words[28]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[28][4] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[6]  ( .D(\words[28]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[28][6] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[8]  ( .D(\words[28]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[28][8] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[10]  ( .D(\words[28]/data_i[10] ), 
        .CLK(clk), .Q(\read_value_mux[28][10] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[12]  ( .D(\words[28]/data_i[12] ), 
        .CLK(clk), .Q(\read_value_mux[28][12] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[20]  ( .D(\words[28]/data_i[20] ), 
        .CLK(clk), .Q(\read_value_mux[28][20] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[3]  ( .D(\words[0]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[0][3] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[5]  ( .D(\words[0]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[0][5] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[7]  ( .D(\words[0]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[0][7] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[9]  ( .D(\words[0]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[0][9] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[11]  ( .D(\words[0]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[0][11] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[13]  ( .D(\words[0]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[0][13] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[15]  ( .D(\words[0]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[0][15] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[17]  ( .D(\words[0]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[0][17] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[19]  ( .D(\words[0]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[0][19] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[21]  ( .D(\words[0]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[0][21] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[23]  ( .D(\words[0]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[0][23] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[25]  ( .D(\words[0]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[0][25] ) );
  DFFX1_RVT \words[0]/data_ff/data_reg[27]  ( .D(\words[0]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[0][27] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[3]  ( .D(\words[3]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[3][3] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[5]  ( .D(\words[3]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[3][5] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[7]  ( .D(\words[3]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[3][7] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[9]  ( .D(\words[3]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[3][9] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[11]  ( .D(\words[3]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[3][11] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[13]  ( .D(\words[3]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[3][13] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[15]  ( .D(\words[3]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[3][15] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[17]  ( .D(\words[3]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[3][17] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[19]  ( .D(\words[3]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[3][19] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[21]  ( .D(\words[3]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[3][21] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[23]  ( .D(\words[3]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[3][23] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[25]  ( .D(\words[3]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[3][25] ) );
  DFFX1_RVT \words[3]/data_ff/data_reg[27]  ( .D(\words[3]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[3][27] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[3]  ( .D(\words[4]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[4][3] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[5]  ( .D(\words[4]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[4][5] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[7]  ( .D(\words[4]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[4][7] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[9]  ( .D(\words[4]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[4][9] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[11]  ( .D(\words[4]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[4][11] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[13]  ( .D(\words[4]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[4][13] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[15]  ( .D(\words[4]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[4][15] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[17]  ( .D(\words[4]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[4][17] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[19]  ( .D(\words[4]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[4][19] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[21]  ( .D(\words[4]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[4][21] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[23]  ( .D(\words[4]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[4][23] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[25]  ( .D(\words[4]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[4][25] ) );
  DFFX1_RVT \words[4]/data_ff/data_reg[27]  ( .D(\words[4]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[4][27] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[3]  ( .D(\words[7]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[7][3] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[5]  ( .D(\words[7]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[7][5] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[7]  ( .D(\words[7]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[7][7] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[11]  ( .D(\words[7]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[7][11] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[13]  ( .D(\words[7]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[7][13] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[15]  ( .D(\words[7]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[7][15] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[19]  ( .D(\words[7]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[7][19] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[21]  ( .D(\words[7]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[7][21] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[27]  ( .D(\words[7]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[7][27] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[3]  ( .D(\words[19]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[19][3] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[5]  ( .D(\words[19]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[19][5] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[7]  ( .D(\words[19]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[19][7] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[9]  ( .D(\words[19]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[19][9] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[11]  ( .D(\words[19]/data_i[11] ), 
        .CLK(clk), .Q(\read_value_mux[19][11] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[13]  ( .D(\words[19]/data_i[13] ), 
        .CLK(clk), .Q(\read_value_mux[19][13] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[15]  ( .D(\words[19]/data_i[15] ), 
        .CLK(clk), .Q(\read_value_mux[19][15] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[17]  ( .D(\words[19]/data_i[17] ), 
        .CLK(clk), .Q(\read_value_mux[19][17] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[19]  ( .D(\words[19]/data_i[19] ), 
        .CLK(clk), .Q(\read_value_mux[19][19] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[21]  ( .D(\words[19]/data_i[21] ), 
        .CLK(clk), .Q(\read_value_mux[19][21] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[23]  ( .D(\words[19]/data_i[23] ), 
        .CLK(clk), .Q(\read_value_mux[19][23] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[25]  ( .D(\words[19]/data_i[25] ), 
        .CLK(clk), .Q(\read_value_mux[19][25] ) );
  DFFX1_RVT \words[19]/data_ff/data_reg[27]  ( .D(\words[19]/data_i[27] ), 
        .CLK(clk), .Q(\read_value_mux[19][27] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[3]  ( .D(\words[28]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[28][3] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[5]  ( .D(\words[28]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[28][5] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[7]  ( .D(\words[28]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[28][7] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[9]  ( .D(\words[28]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[28][9] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[11]  ( .D(\words[28]/data_i[11] ), 
        .CLK(clk), .Q(\read_value_mux[28][11] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[13]  ( .D(\words[28]/data_i[13] ), 
        .CLK(clk), .Q(\read_value_mux[28][13] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[15]  ( .D(\words[28]/data_i[15] ), 
        .CLK(clk), .Q(\read_value_mux[28][15] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[17]  ( .D(\words[28]/data_i[17] ), 
        .CLK(clk), .Q(\read_value_mux[28][17] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[19]  ( .D(\words[28]/data_i[19] ), 
        .CLK(clk), .Q(\read_value_mux[28][19] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[21]  ( .D(\words[28]/data_i[21] ), 
        .CLK(clk), .Q(\read_value_mux[28][21] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[23]  ( .D(\words[28]/data_i[23] ), 
        .CLK(clk), .Q(\read_value_mux[28][23] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[25]  ( .D(\words[28]/data_i[25] ), 
        .CLK(clk), .Q(\read_value_mux[28][25] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[27]  ( .D(\words[28]/data_i[27] ), 
        .CLK(clk), .Q(\read_value_mux[28][27] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[4]  ( .D(\words[5]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[5][4] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[8]  ( .D(\words[5]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[5][8] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[12]  ( .D(\words[5]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[5][12] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[14]  ( .D(\words[5]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[5][14] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[16]  ( .D(\words[5]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[5][16] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[20]  ( .D(\words[5]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[5][20] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[22]  ( .D(\words[5]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[5][22] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[24]  ( .D(\words[5]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[5][24] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[26]  ( .D(\words[5]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[5][26] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[2]  ( .D(\words[10]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[10][2] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[4]  ( .D(\words[10]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[10][4] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[6]  ( .D(\words[10]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[10][6] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[8]  ( .D(\words[10]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[10][8] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[10]  ( .D(\words[10]/data_i[10] ), 
        .CLK(clk), .Q(\read_value_mux[10][10] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[12]  ( .D(\words[10]/data_i[12] ), 
        .CLK(clk), .Q(\read_value_mux[10][12] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[14]  ( .D(\words[10]/data_i[14] ), 
        .CLK(clk), .Q(\read_value_mux[10][14] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[16]  ( .D(\words[10]/data_i[16] ), 
        .CLK(clk), .Q(\read_value_mux[10][16] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[18]  ( .D(\words[10]/data_i[18] ), 
        .CLK(clk), .Q(\read_value_mux[10][18] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[20]  ( .D(\words[10]/data_i[20] ), 
        .CLK(clk), .Q(\read_value_mux[10][20] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[22]  ( .D(\words[10]/data_i[22] ), 
        .CLK(clk), .Q(\read_value_mux[10][22] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[24]  ( .D(\words[10]/data_i[24] ), 
        .CLK(clk), .Q(\read_value_mux[10][24] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[26]  ( .D(\words[10]/data_i[26] ), 
        .CLK(clk), .Q(\read_value_mux[10][26] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[2]  ( .D(\words[13]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[13][2] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[4]  ( .D(\words[13]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[13][4] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[6]  ( .D(\words[13]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[13][6] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[8]  ( .D(\words[13]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[13][8] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[10]  ( .D(\words[13]/data_i[10] ), 
        .CLK(clk), .Q(\read_value_mux[13][10] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[12]  ( .D(\words[13]/data_i[12] ), 
        .CLK(clk), .Q(\read_value_mux[13][12] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[14]  ( .D(\words[13]/data_i[14] ), 
        .CLK(clk), .Q(\read_value_mux[13][14] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[16]  ( .D(\words[13]/data_i[16] ), 
        .CLK(clk), .Q(\read_value_mux[13][16] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[18]  ( .D(\words[13]/data_i[18] ), 
        .CLK(clk), .Q(\read_value_mux[13][18] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[20]  ( .D(\words[13]/data_i[20] ), 
        .CLK(clk), .Q(\read_value_mux[13][20] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[22]  ( .D(\words[13]/data_i[22] ), 
        .CLK(clk), .Q(\read_value_mux[13][22] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[24]  ( .D(\words[13]/data_i[24] ), 
        .CLK(clk), .Q(\read_value_mux[13][24] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[26]  ( .D(\words[13]/data_i[26] ), 
        .CLK(clk), .Q(\read_value_mux[13][26] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[2]  ( .D(\words[14]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[14][2] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[4]  ( .D(\words[14]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[14][4] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[6]  ( .D(\words[14]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[14][6] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[8]  ( .D(\words[14]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[14][8] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[10]  ( .D(\words[14]/data_i[10] ), 
        .CLK(clk), .Q(\read_value_mux[14][10] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[12]  ( .D(\words[14]/data_i[12] ), 
        .CLK(clk), .Q(\read_value_mux[14][12] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[14]  ( .D(\words[14]/data_i[14] ), 
        .CLK(clk), .Q(\read_value_mux[14][14] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[16]  ( .D(\words[14]/data_i[16] ), 
        .CLK(clk), .Q(\read_value_mux[14][16] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[18]  ( .D(\words[14]/data_i[18] ), 
        .CLK(clk), .Q(\read_value_mux[14][18] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[20]  ( .D(\words[14]/data_i[20] ), 
        .CLK(clk), .Q(\read_value_mux[14][20] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[22]  ( .D(\words[14]/data_i[22] ), 
        .CLK(clk), .Q(\read_value_mux[14][22] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[24]  ( .D(\words[14]/data_i[24] ), 
        .CLK(clk), .Q(\read_value_mux[14][24] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[26]  ( .D(\words[14]/data_i[26] ), 
        .CLK(clk), .Q(\read_value_mux[14][26] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[2]  ( .D(\words[18]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[18][2] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[4]  ( .D(\words[18]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[18][4] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[6]  ( .D(\words[18]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[18][6] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[8]  ( .D(\words[18]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[18][8] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[10]  ( .D(\words[18]/data_i[10] ), 
        .CLK(clk), .Q(\read_value_mux[18][10] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[12]  ( .D(\words[18]/data_i[12] ), 
        .CLK(clk), .Q(\read_value_mux[18][12] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[14]  ( .D(\words[18]/data_i[14] ), 
        .CLK(clk), .Q(\read_value_mux[18][14] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[16]  ( .D(\words[18]/data_i[16] ), 
        .CLK(clk), .Q(\read_value_mux[18][16] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[18]  ( .D(\words[18]/data_i[18] ), 
        .CLK(clk), .Q(\read_value_mux[18][18] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[20]  ( .D(\words[18]/data_i[20] ), 
        .CLK(clk), .Q(\read_value_mux[18][20] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[22]  ( .D(\words[18]/data_i[22] ), 
        .CLK(clk), .Q(\read_value_mux[18][22] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[24]  ( .D(\words[18]/data_i[24] ), 
        .CLK(clk), .Q(\read_value_mux[18][24] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[26]  ( .D(\words[18]/data_i[26] ), 
        .CLK(clk), .Q(\read_value_mux[18][26] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[2]  ( .D(\words[21]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[21][2] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[4]  ( .D(\words[21]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[21][4] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[6]  ( .D(\words[21]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[21][6] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[8]  ( .D(\words[21]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[21][8] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[10]  ( .D(\words[21]/data_i[10] ), 
        .CLK(clk), .Q(\read_value_mux[21][10] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[12]  ( .D(\words[21]/data_i[12] ), 
        .CLK(clk), .Q(\read_value_mux[21][12] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[14]  ( .D(\words[21]/data_i[14] ), 
        .CLK(clk), .Q(\read_value_mux[21][14] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[16]  ( .D(\words[21]/data_i[16] ), 
        .CLK(clk), .Q(\read_value_mux[21][16] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[18]  ( .D(\words[21]/data_i[18] ), 
        .CLK(clk), .Q(\read_value_mux[21][18] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[20]  ( .D(\words[21]/data_i[20] ), 
        .CLK(clk), .Q(\read_value_mux[21][20] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[22]  ( .D(\words[21]/data_i[22] ), 
        .CLK(clk), .Q(\read_value_mux[21][22] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[24]  ( .D(\words[21]/data_i[24] ), 
        .CLK(clk), .Q(\read_value_mux[21][24] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[26]  ( .D(\words[21]/data_i[26] ), 
        .CLK(clk), .Q(\read_value_mux[21][26] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[2]  ( .D(\words[22]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[22][2] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[4]  ( .D(\words[22]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[22][4] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[6]  ( .D(\words[22]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[22][6] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[8]  ( .D(\words[22]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[22][8] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[10]  ( .D(\words[22]/data_i[10] ), 
        .CLK(clk), .Q(\read_value_mux[22][10] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[12]  ( .D(\words[22]/data_i[12] ), 
        .CLK(clk), .Q(\read_value_mux[22][12] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[14]  ( .D(\words[22]/data_i[14] ), 
        .CLK(clk), .Q(\read_value_mux[22][14] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[16]  ( .D(\words[22]/data_i[16] ), 
        .CLK(clk), .Q(\read_value_mux[22][16] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[18]  ( .D(\words[22]/data_i[18] ), 
        .CLK(clk), .Q(\read_value_mux[22][18] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[20]  ( .D(\words[22]/data_i[20] ), 
        .CLK(clk), .Q(\read_value_mux[22][20] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[22]  ( .D(\words[22]/data_i[22] ), 
        .CLK(clk), .Q(\read_value_mux[22][22] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[24]  ( .D(\words[22]/data_i[24] ), 
        .CLK(clk), .Q(\read_value_mux[22][24] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[26]  ( .D(\words[22]/data_i[26] ), 
        .CLK(clk), .Q(\read_value_mux[22][26] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[2]  ( .D(\words[25]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[25][2] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[4]  ( .D(\words[25]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[25][4] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[6]  ( .D(\words[25]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[25][6] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[8]  ( .D(\words[25]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[25][8] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[10]  ( .D(\words[25]/data_i[10] ), 
        .CLK(clk), .Q(\read_value_mux[25][10] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[12]  ( .D(\words[25]/data_i[12] ), 
        .CLK(clk), .Q(\read_value_mux[25][12] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[14]  ( .D(\words[25]/data_i[14] ), 
        .CLK(clk), .Q(\read_value_mux[25][14] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[16]  ( .D(\words[25]/data_i[16] ), 
        .CLK(clk), .Q(\read_value_mux[25][16] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[18]  ( .D(\words[25]/data_i[18] ), 
        .CLK(clk), .Q(\read_value_mux[25][18] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[20]  ( .D(\words[25]/data_i[20] ), 
        .CLK(clk), .Q(\read_value_mux[25][20] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[22]  ( .D(\words[25]/data_i[22] ), 
        .CLK(clk), .Q(\read_value_mux[25][22] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[24]  ( .D(\words[25]/data_i[24] ), 
        .CLK(clk), .Q(\read_value_mux[25][24] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[26]  ( .D(\words[25]/data_i[26] ), 
        .CLK(clk), .Q(\read_value_mux[25][26] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[2]  ( .D(\words[26]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[26][2] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[4]  ( .D(\words[26]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[26][4] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[6]  ( .D(\words[26]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[26][6] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[8]  ( .D(\words[26]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[26][8] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[10]  ( .D(\words[26]/data_i[10] ), 
        .CLK(clk), .Q(\read_value_mux[26][10] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[12]  ( .D(\words[26]/data_i[12] ), 
        .CLK(clk), .Q(\read_value_mux[26][12] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[14]  ( .D(\words[26]/data_i[14] ), 
        .CLK(clk), .Q(\read_value_mux[26][14] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[16]  ( .D(\words[26]/data_i[16] ), 
        .CLK(clk), .Q(\read_value_mux[26][16] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[18]  ( .D(\words[26]/data_i[18] ), 
        .CLK(clk), .Q(\read_value_mux[26][18] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[20]  ( .D(\words[26]/data_i[20] ), 
        .CLK(clk), .Q(\read_value_mux[26][20] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[22]  ( .D(\words[26]/data_i[22] ), 
        .CLK(clk), .Q(\read_value_mux[26][22] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[24]  ( .D(\words[26]/data_i[24] ), 
        .CLK(clk), .Q(\read_value_mux[26][24] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[26]  ( .D(\words[26]/data_i[26] ), 
        .CLK(clk), .Q(\read_value_mux[26][26] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[2]  ( .D(\words[29]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[29][2] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[4]  ( .D(\words[29]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[29][4] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[6]  ( .D(\words[29]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[29][6] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[8]  ( .D(\words[29]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[29][8] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[10]  ( .D(\words[29]/data_i[10] ), 
        .CLK(clk), .Q(\read_value_mux[29][10] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[12]  ( .D(\words[29]/data_i[12] ), 
        .CLK(clk), .Q(\read_value_mux[29][12] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[14]  ( .D(\words[29]/data_i[14] ), 
        .CLK(clk), .Q(\read_value_mux[29][14] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[16]  ( .D(\words[29]/data_i[16] ), 
        .CLK(clk), .Q(\read_value_mux[29][16] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[18]  ( .D(\words[29]/data_i[18] ), 
        .CLK(clk), .Q(\read_value_mux[29][18] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[20]  ( .D(\words[29]/data_i[20] ), 
        .CLK(clk), .Q(\read_value_mux[29][20] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[22]  ( .D(\words[29]/data_i[22] ), 
        .CLK(clk), .Q(\read_value_mux[29][22] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[24]  ( .D(\words[29]/data_i[24] ), 
        .CLK(clk), .Q(\read_value_mux[29][24] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[26]  ( .D(\words[29]/data_i[26] ), 
        .CLK(clk), .Q(\read_value_mux[29][26] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[2]  ( .D(\words[30]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[30][2] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[4]  ( .D(\words[30]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[30][4] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[6]  ( .D(\words[30]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[30][6] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[8]  ( .D(\words[30]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[30][8] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[10]  ( .D(\words[30]/data_i[10] ), 
        .CLK(clk), .Q(\read_value_mux[30][10] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[12]  ( .D(\words[30]/data_i[12] ), 
        .CLK(clk), .Q(\read_value_mux[30][12] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[14]  ( .D(\words[30]/data_i[14] ), 
        .CLK(clk), .Q(\read_value_mux[30][14] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[16]  ( .D(\words[30]/data_i[16] ), 
        .CLK(clk), .Q(\read_value_mux[30][16] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[18]  ( .D(\words[30]/data_i[18] ), 
        .CLK(clk), .Q(\read_value_mux[30][18] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[20]  ( .D(\words[30]/data_i[20] ), 
        .CLK(clk), .Q(\read_value_mux[30][20] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[22]  ( .D(\words[30]/data_i[22] ), 
        .CLK(clk), .Q(\read_value_mux[30][22] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[24]  ( .D(\words[30]/data_i[24] ), 
        .CLK(clk), .Q(\read_value_mux[30][24] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[26]  ( .D(\words[30]/data_i[26] ), 
        .CLK(clk), .Q(\read_value_mux[30][26] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[0]  ( .D(\words[9]/data_i[0] ), .CLK(
        clk), .Q(\read_value_mux[9][0] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[1]  ( .D(\words[9]/data_i[1] ), .CLK(
        clk), .Q(\read_value_mux[9][1] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[2]  ( .D(\words[9]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[9][2] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[4]  ( .D(\words[9]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[9][4] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[6]  ( .D(\words[9]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[9][6] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[8]  ( .D(\words[9]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[9][8] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[10]  ( .D(\words[9]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[9][10] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[12]  ( .D(\words[9]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[9][12] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[14]  ( .D(\words[9]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[9][14] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[16]  ( .D(\words[9]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[9][16] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[18]  ( .D(\words[9]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[9][18] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[20]  ( .D(\words[9]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[9][20] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[22]  ( .D(\words[9]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[9][22] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[24]  ( .D(\words[9]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[9][24] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[26]  ( .D(\words[9]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[9][26] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[3]  ( .D(\words[9]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[9][3] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[5]  ( .D(\words[9]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[9][5] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[7]  ( .D(\words[9]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[9][7] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[9]  ( .D(\words[9]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[9][9] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[11]  ( .D(\words[9]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[9][11] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[13]  ( .D(\words[9]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[9][13] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[15]  ( .D(\words[9]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[9][15] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[17]  ( .D(\words[9]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[9][17] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[19]  ( .D(\words[9]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[9][19] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[21]  ( .D(\words[9]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[9][21] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[23]  ( .D(\words[9]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[9][23] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[25]  ( .D(\words[9]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[9][25] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[27]  ( .D(\words[9]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[9][27] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[29]  ( .D(\words[9]/data_i[29] ), .CLK(
        clk), .Q(\read_value_mux[9][29] ) );
  DFFX1_RVT \words[9]/data_ff/data_reg[31]  ( .D(\words[9]/data_i[31] ), .CLK(
        clk), .Q(\read_value_mux[9][31] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[5]  ( .D(\words[5]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[5][5] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[9]  ( .D(\words[5]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[5][9] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[13]  ( .D(\words[5]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[5][13] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[15]  ( .D(\words[5]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[5][15] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[17]  ( .D(\words[5]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[5][17] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[21]  ( .D(\words[5]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[5][21] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[23]  ( .D(\words[5]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[5][23] ) );
  DFFX1_RVT \words[5]/data_ff/data_reg[25]  ( .D(\words[5]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[5][25] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[3]  ( .D(\words[10]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[10][3] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[7]  ( .D(\words[10]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[10][7] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[9]  ( .D(\words[10]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[10][9] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[11]  ( .D(\words[10]/data_i[11] ), 
        .CLK(clk), .Q(\read_value_mux[10][11] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[15]  ( .D(\words[10]/data_i[15] ), 
        .CLK(clk), .Q(\read_value_mux[10][15] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[17]  ( .D(\words[10]/data_i[17] ), 
        .CLK(clk), .Q(\read_value_mux[10][17] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[19]  ( .D(\words[10]/data_i[19] ), 
        .CLK(clk), .Q(\read_value_mux[10][19] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[21]  ( .D(\words[10]/data_i[21] ), 
        .CLK(clk), .Q(\read_value_mux[10][21] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[23]  ( .D(\words[10]/data_i[23] ), 
        .CLK(clk), .Q(\read_value_mux[10][23] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[25]  ( .D(\words[10]/data_i[25] ), 
        .CLK(clk), .Q(\read_value_mux[10][25] ) );
  DFFX1_RVT \words[10]/data_ff/data_reg[27]  ( .D(\words[10]/data_i[27] ), 
        .CLK(clk), .Q(\read_value_mux[10][27] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[3]  ( .D(\words[13]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[13][3] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[5]  ( .D(\words[13]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[13][5] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[7]  ( .D(\words[13]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[13][7] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[9]  ( .D(\words[13]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[13][9] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[11]  ( .D(\words[13]/data_i[11] ), 
        .CLK(clk), .Q(\read_value_mux[13][11] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[13]  ( .D(\words[13]/data_i[13] ), 
        .CLK(clk), .Q(\read_value_mux[13][13] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[15]  ( .D(\words[13]/data_i[15] ), 
        .CLK(clk), .Q(\read_value_mux[13][15] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[17]  ( .D(\words[13]/data_i[17] ), 
        .CLK(clk), .Q(\read_value_mux[13][17] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[19]  ( .D(\words[13]/data_i[19] ), 
        .CLK(clk), .Q(\read_value_mux[13][19] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[21]  ( .D(\words[13]/data_i[21] ), 
        .CLK(clk), .Q(\read_value_mux[13][21] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[23]  ( .D(\words[13]/data_i[23] ), 
        .CLK(clk), .Q(\read_value_mux[13][23] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[25]  ( .D(\words[13]/data_i[25] ), 
        .CLK(clk), .Q(\read_value_mux[13][25] ) );
  DFFX1_RVT \words[13]/data_ff/data_reg[27]  ( .D(\words[13]/data_i[27] ), 
        .CLK(clk), .Q(\read_value_mux[13][27] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[3]  ( .D(\words[14]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[14][3] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[5]  ( .D(\words[14]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[14][5] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[7]  ( .D(\words[14]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[14][7] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[9]  ( .D(\words[14]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[14][9] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[11]  ( .D(\words[14]/data_i[11] ), 
        .CLK(clk), .Q(\read_value_mux[14][11] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[13]  ( .D(\words[14]/data_i[13] ), 
        .CLK(clk), .Q(\read_value_mux[14][13] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[15]  ( .D(\words[14]/data_i[15] ), 
        .CLK(clk), .Q(\read_value_mux[14][15] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[17]  ( .D(\words[14]/data_i[17] ), 
        .CLK(clk), .Q(\read_value_mux[14][17] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[19]  ( .D(\words[14]/data_i[19] ), 
        .CLK(clk), .Q(\read_value_mux[14][19] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[21]  ( .D(\words[14]/data_i[21] ), 
        .CLK(clk), .Q(\read_value_mux[14][21] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[23]  ( .D(\words[14]/data_i[23] ), 
        .CLK(clk), .Q(\read_value_mux[14][23] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[25]  ( .D(\words[14]/data_i[25] ), 
        .CLK(clk), .Q(\read_value_mux[14][25] ) );
  DFFX1_RVT \words[14]/data_ff/data_reg[27]  ( .D(\words[14]/data_i[27] ), 
        .CLK(clk), .Q(\read_value_mux[14][27] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[3]  ( .D(\words[18]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[18][3] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[5]  ( .D(\words[18]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[18][5] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[7]  ( .D(\words[18]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[18][7] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[9]  ( .D(\words[18]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[18][9] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[11]  ( .D(\words[18]/data_i[11] ), 
        .CLK(clk), .Q(\read_value_mux[18][11] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[13]  ( .D(\words[18]/data_i[13] ), 
        .CLK(clk), .Q(\read_value_mux[18][13] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[15]  ( .D(\words[18]/data_i[15] ), 
        .CLK(clk), .Q(\read_value_mux[18][15] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[17]  ( .D(\words[18]/data_i[17] ), 
        .CLK(clk), .Q(\read_value_mux[18][17] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[19]  ( .D(\words[18]/data_i[19] ), 
        .CLK(clk), .Q(\read_value_mux[18][19] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[21]  ( .D(\words[18]/data_i[21] ), 
        .CLK(clk), .Q(\read_value_mux[18][21] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[23]  ( .D(\words[18]/data_i[23] ), 
        .CLK(clk), .Q(\read_value_mux[18][23] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[25]  ( .D(\words[18]/data_i[25] ), 
        .CLK(clk), .Q(\read_value_mux[18][25] ) );
  DFFX1_RVT \words[18]/data_ff/data_reg[27]  ( .D(\words[18]/data_i[27] ), 
        .CLK(clk), .Q(\read_value_mux[18][27] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[3]  ( .D(\words[21]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[21][3] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[5]  ( .D(\words[21]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[21][5] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[7]  ( .D(\words[21]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[21][7] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[9]  ( .D(\words[21]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[21][9] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[11]  ( .D(\words[21]/data_i[11] ), 
        .CLK(clk), .Q(\read_value_mux[21][11] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[13]  ( .D(\words[21]/data_i[13] ), 
        .CLK(clk), .Q(\read_value_mux[21][13] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[15]  ( .D(\words[21]/data_i[15] ), 
        .CLK(clk), .Q(\read_value_mux[21][15] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[17]  ( .D(\words[21]/data_i[17] ), 
        .CLK(clk), .Q(\read_value_mux[21][17] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[19]  ( .D(\words[21]/data_i[19] ), 
        .CLK(clk), .Q(\read_value_mux[21][19] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[21]  ( .D(\words[21]/data_i[21] ), 
        .CLK(clk), .Q(\read_value_mux[21][21] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[23]  ( .D(\words[21]/data_i[23] ), 
        .CLK(clk), .Q(\read_value_mux[21][23] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[25]  ( .D(\words[21]/data_i[25] ), 
        .CLK(clk), .Q(\read_value_mux[21][25] ) );
  DFFX1_RVT \words[21]/data_ff/data_reg[27]  ( .D(\words[21]/data_i[27] ), 
        .CLK(clk), .Q(\read_value_mux[21][27] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[3]  ( .D(\words[22]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[22][3] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[5]  ( .D(\words[22]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[22][5] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[7]  ( .D(\words[22]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[22][7] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[9]  ( .D(\words[22]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[22][9] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[11]  ( .D(\words[22]/data_i[11] ), 
        .CLK(clk), .Q(\read_value_mux[22][11] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[13]  ( .D(\words[22]/data_i[13] ), 
        .CLK(clk), .Q(\read_value_mux[22][13] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[15]  ( .D(\words[22]/data_i[15] ), 
        .CLK(clk), .Q(\read_value_mux[22][15] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[17]  ( .D(\words[22]/data_i[17] ), 
        .CLK(clk), .Q(\read_value_mux[22][17] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[19]  ( .D(\words[22]/data_i[19] ), 
        .CLK(clk), .Q(\read_value_mux[22][19] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[21]  ( .D(\words[22]/data_i[21] ), 
        .CLK(clk), .Q(\read_value_mux[22][21] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[23]  ( .D(\words[22]/data_i[23] ), 
        .CLK(clk), .Q(\read_value_mux[22][23] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[25]  ( .D(\words[22]/data_i[25] ), 
        .CLK(clk), .Q(\read_value_mux[22][25] ) );
  DFFX1_RVT \words[22]/data_ff/data_reg[27]  ( .D(\words[22]/data_i[27] ), 
        .CLK(clk), .Q(\read_value_mux[22][27] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[3]  ( .D(\words[25]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[25][3] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[5]  ( .D(\words[25]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[25][5] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[7]  ( .D(\words[25]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[25][7] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[9]  ( .D(\words[25]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[25][9] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[11]  ( .D(\words[25]/data_i[11] ), 
        .CLK(clk), .Q(\read_value_mux[25][11] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[13]  ( .D(\words[25]/data_i[13] ), 
        .CLK(clk), .Q(\read_value_mux[25][13] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[15]  ( .D(\words[25]/data_i[15] ), 
        .CLK(clk), .Q(\read_value_mux[25][15] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[17]  ( .D(\words[25]/data_i[17] ), 
        .CLK(clk), .Q(\read_value_mux[25][17] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[19]  ( .D(\words[25]/data_i[19] ), 
        .CLK(clk), .Q(\read_value_mux[25][19] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[21]  ( .D(\words[25]/data_i[21] ), 
        .CLK(clk), .Q(\read_value_mux[25][21] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[23]  ( .D(\words[25]/data_i[23] ), 
        .CLK(clk), .Q(\read_value_mux[25][23] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[25]  ( .D(\words[25]/data_i[25] ), 
        .CLK(clk), .Q(\read_value_mux[25][25] ) );
  DFFX1_RVT \words[25]/data_ff/data_reg[27]  ( .D(\words[25]/data_i[27] ), 
        .CLK(clk), .Q(\read_value_mux[25][27] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[3]  ( .D(\words[26]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[26][3] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[5]  ( .D(\words[26]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[26][5] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[7]  ( .D(\words[26]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[26][7] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[9]  ( .D(\words[26]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[26][9] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[11]  ( .D(\words[26]/data_i[11] ), 
        .CLK(clk), .Q(\read_value_mux[26][11] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[13]  ( .D(\words[26]/data_i[13] ), 
        .CLK(clk), .Q(\read_value_mux[26][13] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[15]  ( .D(\words[26]/data_i[15] ), 
        .CLK(clk), .Q(\read_value_mux[26][15] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[17]  ( .D(\words[26]/data_i[17] ), 
        .CLK(clk), .Q(\read_value_mux[26][17] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[19]  ( .D(\words[26]/data_i[19] ), 
        .CLK(clk), .Q(\read_value_mux[26][19] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[21]  ( .D(\words[26]/data_i[21] ), 
        .CLK(clk), .Q(\read_value_mux[26][21] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[23]  ( .D(\words[26]/data_i[23] ), 
        .CLK(clk), .Q(\read_value_mux[26][23] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[25]  ( .D(\words[26]/data_i[25] ), 
        .CLK(clk), .Q(\read_value_mux[26][25] ) );
  DFFX1_RVT \words[26]/data_ff/data_reg[27]  ( .D(\words[26]/data_i[27] ), 
        .CLK(clk), .Q(\read_value_mux[26][27] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[3]  ( .D(\words[29]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[29][3] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[5]  ( .D(\words[29]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[29][5] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[7]  ( .D(\words[29]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[29][7] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[9]  ( .D(\words[29]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[29][9] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[11]  ( .D(\words[29]/data_i[11] ), 
        .CLK(clk), .Q(\read_value_mux[29][11] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[13]  ( .D(\words[29]/data_i[13] ), 
        .CLK(clk), .Q(\read_value_mux[29][13] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[15]  ( .D(\words[29]/data_i[15] ), 
        .CLK(clk), .Q(\read_value_mux[29][15] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[17]  ( .D(\words[29]/data_i[17] ), 
        .CLK(clk), .Q(\read_value_mux[29][17] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[19]  ( .D(\words[29]/data_i[19] ), 
        .CLK(clk), .Q(\read_value_mux[29][19] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[21]  ( .D(\words[29]/data_i[21] ), 
        .CLK(clk), .Q(\read_value_mux[29][21] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[23]  ( .D(\words[29]/data_i[23] ), 
        .CLK(clk), .Q(\read_value_mux[29][23] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[25]  ( .D(\words[29]/data_i[25] ), 
        .CLK(clk), .Q(\read_value_mux[29][25] ) );
  DFFX1_RVT \words[29]/data_ff/data_reg[27]  ( .D(\words[29]/data_i[27] ), 
        .CLK(clk), .Q(\read_value_mux[29][27] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[3]  ( .D(\words[30]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[30][3] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[5]  ( .D(\words[30]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[30][5] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[7]  ( .D(\words[30]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[30][7] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[9]  ( .D(\words[30]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[30][9] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[11]  ( .D(\words[30]/data_i[11] ), 
        .CLK(clk), .Q(\read_value_mux[30][11] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[13]  ( .D(\words[30]/data_i[13] ), 
        .CLK(clk), .Q(\read_value_mux[30][13] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[15]  ( .D(\words[30]/data_i[15] ), 
        .CLK(clk), .Q(\read_value_mux[30][15] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[17]  ( .D(\words[30]/data_i[17] ), 
        .CLK(clk), .Q(\read_value_mux[30][17] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[19]  ( .D(\words[30]/data_i[19] ), 
        .CLK(clk), .Q(\read_value_mux[30][19] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[21]  ( .D(\words[30]/data_i[21] ), 
        .CLK(clk), .Q(\read_value_mux[30][21] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[23]  ( .D(\words[30]/data_i[23] ), 
        .CLK(clk), .Q(\read_value_mux[30][23] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[25]  ( .D(\words[30]/data_i[25] ), 
        .CLK(clk), .Q(\read_value_mux[30][25] ) );
  DFFX1_RVT \words[30]/data_ff/data_reg[27]  ( .D(\words[30]/data_i[27] ), 
        .CLK(clk), .Q(\read_value_mux[30][27] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[2]  ( .D(\words[31]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[31][2] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[4]  ( .D(\words[31]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[31][4] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[6]  ( .D(\words[31]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[31][6] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[8]  ( .D(\words[31]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[31][8] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[10]  ( .D(\words[31]/data_i[10] ), 
        .CLK(clk), .Q(\read_value_mux[31][10] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[12]  ( .D(\words[31]/data_i[12] ), 
        .CLK(clk), .Q(\read_value_mux[31][12] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[14]  ( .D(\words[31]/data_i[14] ), 
        .CLK(clk), .Q(\read_value_mux[31][14] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[16]  ( .D(\words[31]/data_i[16] ), 
        .CLK(clk), .Q(\read_value_mux[31][16] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[18]  ( .D(\words[31]/data_i[18] ), 
        .CLK(clk), .Q(\read_value_mux[31][18] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[20]  ( .D(\words[31]/data_i[20] ), 
        .CLK(clk), .Q(\read_value_mux[31][20] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[22]  ( .D(\words[31]/data_i[22] ), 
        .CLK(clk), .Q(\read_value_mux[31][22] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[24]  ( .D(\words[31]/data_i[24] ), 
        .CLK(clk), .Q(\read_value_mux[31][24] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[26]  ( .D(\words[31]/data_i[26] ), 
        .CLK(clk), .Q(\read_value_mux[31][26] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[4]  ( .D(\words[7]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[7][4] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[8]  ( .D(\words[7]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[7][8] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[12]  ( .D(\words[7]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[7][12] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[14]  ( .D(\words[7]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[7][14] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[16]  ( .D(\words[7]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[7][16] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[20]  ( .D(\words[7]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[7][20] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[22]  ( .D(\words[7]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[7][22] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[24]  ( .D(\words[7]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[7][24] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[2]  ( .D(\words[8]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[8][2] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[4]  ( .D(\words[8]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[8][4] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[6]  ( .D(\words[8]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[8][6] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[8]  ( .D(\words[8]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[8][8] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[10]  ( .D(\words[8]/data_i[10] ), .CLK(
        clk), .Q(\read_value_mux[8][10] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[12]  ( .D(\words[8]/data_i[12] ), .CLK(
        clk), .Q(\read_value_mux[8][12] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[14]  ( .D(\words[8]/data_i[14] ), .CLK(
        clk), .Q(\read_value_mux[8][14] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[16]  ( .D(\words[8]/data_i[16] ), .CLK(
        clk), .Q(\read_value_mux[8][16] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[18]  ( .D(\words[8]/data_i[18] ), .CLK(
        clk), .Q(\read_value_mux[8][18] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[20]  ( .D(\words[8]/data_i[20] ), .CLK(
        clk), .Q(\read_value_mux[8][20] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[22]  ( .D(\words[8]/data_i[22] ), .CLK(
        clk), .Q(\read_value_mux[8][22] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[24]  ( .D(\words[8]/data_i[24] ), .CLK(
        clk), .Q(\read_value_mux[8][24] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[26]  ( .D(\words[8]/data_i[26] ), .CLK(
        clk), .Q(\read_value_mux[8][26] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[2]  ( .D(\words[11]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[11][2] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[4]  ( .D(\words[11]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[11][4] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[6]  ( .D(\words[11]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[11][6] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[8]  ( .D(\words[11]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[11][8] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[10]  ( .D(\words[11]/data_i[10] ), 
        .CLK(clk), .Q(\read_value_mux[11][10] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[12]  ( .D(\words[11]/data_i[12] ), 
        .CLK(clk), .Q(\read_value_mux[11][12] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[14]  ( .D(\words[11]/data_i[14] ), 
        .CLK(clk), .Q(\read_value_mux[11][14] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[16]  ( .D(\words[11]/data_i[16] ), 
        .CLK(clk), .Q(\read_value_mux[11][16] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[18]  ( .D(\words[11]/data_i[18] ), 
        .CLK(clk), .Q(\read_value_mux[11][18] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[20]  ( .D(\words[11]/data_i[20] ), 
        .CLK(clk), .Q(\read_value_mux[11][20] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[22]  ( .D(\words[11]/data_i[22] ), 
        .CLK(clk), .Q(\read_value_mux[11][22] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[24]  ( .D(\words[11]/data_i[24] ), 
        .CLK(clk), .Q(\read_value_mux[11][24] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[26]  ( .D(\words[11]/data_i[26] ), 
        .CLK(clk), .Q(\read_value_mux[11][26] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[2]  ( .D(\words[12]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[12][2] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[4]  ( .D(\words[12]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[12][4] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[6]  ( .D(\words[12]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[12][6] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[8]  ( .D(\words[12]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[12][8] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[10]  ( .D(\words[12]/data_i[10] ), 
        .CLK(clk), .Q(\read_value_mux[12][10] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[12]  ( .D(\words[12]/data_i[12] ), 
        .CLK(clk), .Q(\read_value_mux[12][12] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[14]  ( .D(\words[12]/data_i[14] ), 
        .CLK(clk), .Q(\read_value_mux[12][14] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[16]  ( .D(\words[12]/data_i[16] ), 
        .CLK(clk), .Q(\read_value_mux[12][16] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[18]  ( .D(\words[12]/data_i[18] ), 
        .CLK(clk), .Q(\read_value_mux[12][18] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[20]  ( .D(\words[12]/data_i[20] ), 
        .CLK(clk), .Q(\read_value_mux[12][20] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[22]  ( .D(\words[12]/data_i[22] ), 
        .CLK(clk), .Q(\read_value_mux[12][22] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[24]  ( .D(\words[12]/data_i[24] ), 
        .CLK(clk), .Q(\read_value_mux[12][24] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[26]  ( .D(\words[12]/data_i[26] ), 
        .CLK(clk), .Q(\read_value_mux[12][26] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[2]  ( .D(\words[15]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[15][2] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[4]  ( .D(\words[15]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[15][4] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[6]  ( .D(\words[15]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[15][6] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[8]  ( .D(\words[15]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[15][8] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[10]  ( .D(\words[15]/data_i[10] ), 
        .CLK(clk), .Q(\read_value_mux[15][10] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[12]  ( .D(\words[15]/data_i[12] ), 
        .CLK(clk), .Q(\read_value_mux[15][12] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[14]  ( .D(\words[15]/data_i[14] ), 
        .CLK(clk), .Q(\read_value_mux[15][14] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[16]  ( .D(\words[15]/data_i[16] ), 
        .CLK(clk), .Q(\read_value_mux[15][16] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[18]  ( .D(\words[15]/data_i[18] ), 
        .CLK(clk), .Q(\read_value_mux[15][18] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[20]  ( .D(\words[15]/data_i[20] ), 
        .CLK(clk), .Q(\read_value_mux[15][20] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[22]  ( .D(\words[15]/data_i[22] ), 
        .CLK(clk), .Q(\read_value_mux[15][22] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[24]  ( .D(\words[15]/data_i[24] ), 
        .CLK(clk), .Q(\read_value_mux[15][24] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[26]  ( .D(\words[15]/data_i[26] ), 
        .CLK(clk), .Q(\read_value_mux[15][26] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[2]  ( .D(\words[16]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[16][2] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[4]  ( .D(\words[16]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[16][4] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[6]  ( .D(\words[16]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[16][6] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[8]  ( .D(\words[16]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[16][8] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[10]  ( .D(\words[16]/data_i[10] ), 
        .CLK(clk), .Q(\read_value_mux[16][10] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[12]  ( .D(\words[16]/data_i[12] ), 
        .CLK(clk), .Q(\read_value_mux[16][12] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[14]  ( .D(\words[16]/data_i[14] ), 
        .CLK(clk), .Q(\read_value_mux[16][14] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[16]  ( .D(\words[16]/data_i[16] ), 
        .CLK(clk), .Q(\read_value_mux[16][16] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[18]  ( .D(\words[16]/data_i[18] ), 
        .CLK(clk), .Q(\read_value_mux[16][18] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[20]  ( .D(\words[16]/data_i[20] ), 
        .CLK(clk), .Q(\read_value_mux[16][20] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[22]  ( .D(\words[16]/data_i[22] ), 
        .CLK(clk), .Q(\read_value_mux[16][22] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[24]  ( .D(\words[16]/data_i[24] ), 
        .CLK(clk), .Q(\read_value_mux[16][24] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[26]  ( .D(\words[16]/data_i[26] ), 
        .CLK(clk), .Q(\read_value_mux[16][26] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[2]  ( .D(\words[20]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[20][2] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[4]  ( .D(\words[20]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[20][4] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[6]  ( .D(\words[20]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[20][6] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[8]  ( .D(\words[20]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[20][8] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[10]  ( .D(\words[20]/data_i[10] ), 
        .CLK(clk), .Q(\read_value_mux[20][10] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[12]  ( .D(\words[20]/data_i[12] ), 
        .CLK(clk), .Q(\read_value_mux[20][12] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[14]  ( .D(\words[20]/data_i[14] ), 
        .CLK(clk), .Q(\read_value_mux[20][14] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[16]  ( .D(\words[20]/data_i[16] ), 
        .CLK(clk), .Q(\read_value_mux[20][16] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[18]  ( .D(\words[20]/data_i[18] ), 
        .CLK(clk), .Q(\read_value_mux[20][18] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[20]  ( .D(\words[20]/data_i[20] ), 
        .CLK(clk), .Q(\read_value_mux[20][20] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[22]  ( .D(\words[20]/data_i[22] ), 
        .CLK(clk), .Q(\read_value_mux[20][22] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[24]  ( .D(\words[20]/data_i[24] ), 
        .CLK(clk), .Q(\read_value_mux[20][24] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[26]  ( .D(\words[20]/data_i[26] ), 
        .CLK(clk), .Q(\read_value_mux[20][26] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[2]  ( .D(\words[23]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[23][2] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[4]  ( .D(\words[23]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[23][4] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[6]  ( .D(\words[23]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[23][6] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[8]  ( .D(\words[23]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[23][8] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[10]  ( .D(\words[23]/data_i[10] ), 
        .CLK(clk), .Q(\read_value_mux[23][10] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[12]  ( .D(\words[23]/data_i[12] ), 
        .CLK(clk), .Q(\read_value_mux[23][12] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[14]  ( .D(\words[23]/data_i[14] ), 
        .CLK(clk), .Q(\read_value_mux[23][14] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[16]  ( .D(\words[23]/data_i[16] ), 
        .CLK(clk), .Q(\read_value_mux[23][16] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[18]  ( .D(\words[23]/data_i[18] ), 
        .CLK(clk), .Q(\read_value_mux[23][18] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[20]  ( .D(\words[23]/data_i[20] ), 
        .CLK(clk), .Q(\read_value_mux[23][20] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[22]  ( .D(\words[23]/data_i[22] ), 
        .CLK(clk), .Q(\read_value_mux[23][22] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[24]  ( .D(\words[23]/data_i[24] ), 
        .CLK(clk), .Q(\read_value_mux[23][24] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[26]  ( .D(\words[23]/data_i[26] ), 
        .CLK(clk), .Q(\read_value_mux[23][26] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[2]  ( .D(\words[24]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[24][2] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[4]  ( .D(\words[24]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[24][4] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[6]  ( .D(\words[24]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[24][6] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[8]  ( .D(\words[24]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[24][8] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[10]  ( .D(\words[24]/data_i[10] ), 
        .CLK(clk), .Q(\read_value_mux[24][10] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[12]  ( .D(\words[24]/data_i[12] ), 
        .CLK(clk), .Q(\read_value_mux[24][12] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[14]  ( .D(\words[24]/data_i[14] ), 
        .CLK(clk), .Q(\read_value_mux[24][14] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[16]  ( .D(\words[24]/data_i[16] ), 
        .CLK(clk), .Q(\read_value_mux[24][16] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[18]  ( .D(\words[24]/data_i[18] ), 
        .CLK(clk), .Q(\read_value_mux[24][18] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[20]  ( .D(\words[24]/data_i[20] ), 
        .CLK(clk), .Q(\read_value_mux[24][20] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[22]  ( .D(\words[24]/data_i[22] ), 
        .CLK(clk), .Q(\read_value_mux[24][22] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[24]  ( .D(\words[24]/data_i[24] ), 
        .CLK(clk), .Q(\read_value_mux[24][24] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[26]  ( .D(\words[24]/data_i[26] ), 
        .CLK(clk), .Q(\read_value_mux[24][26] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[2]  ( .D(\words[27]/data_i[2] ), .CLK(
        clk), .Q(\read_value_mux[27][2] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[4]  ( .D(\words[27]/data_i[4] ), .CLK(
        clk), .Q(\read_value_mux[27][4] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[6]  ( .D(\words[27]/data_i[6] ), .CLK(
        clk), .Q(\read_value_mux[27][6] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[8]  ( .D(\words[27]/data_i[8] ), .CLK(
        clk), .Q(\read_value_mux[27][8] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[10]  ( .D(\words[27]/data_i[10] ), 
        .CLK(clk), .Q(\read_value_mux[27][10] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[12]  ( .D(\words[27]/data_i[12] ), 
        .CLK(clk), .Q(\read_value_mux[27][12] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[14]  ( .D(\words[27]/data_i[14] ), 
        .CLK(clk), .Q(\read_value_mux[27][14] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[16]  ( .D(\words[27]/data_i[16] ), 
        .CLK(clk), .Q(\read_value_mux[27][16] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[18]  ( .D(\words[27]/data_i[18] ), 
        .CLK(clk), .Q(\read_value_mux[27][18] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[20]  ( .D(\words[27]/data_i[20] ), 
        .CLK(clk), .Q(\read_value_mux[27][20] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[22]  ( .D(\words[27]/data_i[22] ), 
        .CLK(clk), .Q(\read_value_mux[27][22] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[24]  ( .D(\words[27]/data_i[24] ), 
        .CLK(clk), .Q(\read_value_mux[27][24] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[26]  ( .D(\words[27]/data_i[26] ), 
        .CLK(clk), .Q(\read_value_mux[27][26] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[14]  ( .D(\words[28]/data_i[14] ), 
        .CLK(clk), .Q(\read_value_mux[28][14] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[16]  ( .D(\words[28]/data_i[16] ), 
        .CLK(clk), .Q(\read_value_mux[28][16] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[18]  ( .D(\words[28]/data_i[18] ), 
        .CLK(clk), .Q(\read_value_mux[28][18] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[22]  ( .D(\words[28]/data_i[22] ), 
        .CLK(clk), .Q(\read_value_mux[28][22] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[24]  ( .D(\words[28]/data_i[24] ), 
        .CLK(clk), .Q(\read_value_mux[28][24] ) );
  DFFX1_RVT \words[28]/data_ff/data_reg[26]  ( .D(\words[28]/data_i[26] ), 
        .CLK(clk), .Q(\read_value_mux[28][26] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[3]  ( .D(\words[31]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[31][3] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[5]  ( .D(\words[31]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[31][5] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[7]  ( .D(\words[31]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[31][7] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[9]  ( .D(\words[31]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[31][9] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[11]  ( .D(\words[31]/data_i[11] ), 
        .CLK(clk), .Q(\read_value_mux[31][11] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[13]  ( .D(\words[31]/data_i[13] ), 
        .CLK(clk), .Q(\read_value_mux[31][13] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[15]  ( .D(\words[31]/data_i[15] ), 
        .CLK(clk), .Q(\read_value_mux[31][15] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[17]  ( .D(\words[31]/data_i[17] ), 
        .CLK(clk), .Q(\read_value_mux[31][17] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[19]  ( .D(\words[31]/data_i[19] ), 
        .CLK(clk), .Q(\read_value_mux[31][19] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[21]  ( .D(\words[31]/data_i[21] ), 
        .CLK(clk), .Q(\read_value_mux[31][21] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[23]  ( .D(\words[31]/data_i[23] ), 
        .CLK(clk), .Q(\read_value_mux[31][23] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[25]  ( .D(\words[31]/data_i[25] ), 
        .CLK(clk), .Q(\read_value_mux[31][25] ) );
  DFFX1_RVT \words[31]/data_ff/data_reg[27]  ( .D(\words[31]/data_i[27] ), 
        .CLK(clk), .Q(\read_value_mux[31][27] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[9]  ( .D(\words[7]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[7][9] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[17]  ( .D(\words[7]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[7][17] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[23]  ( .D(\words[7]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[7][23] ) );
  DFFX1_RVT \words[7]/data_ff/data_reg[25]  ( .D(\words[7]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[7][25] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[3]  ( .D(\words[8]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[8][3] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[5]  ( .D(\words[8]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[8][5] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[7]  ( .D(\words[8]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[8][7] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[9]  ( .D(\words[8]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[8][9] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[11]  ( .D(\words[8]/data_i[11] ), .CLK(
        clk), .Q(\read_value_mux[8][11] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[13]  ( .D(\words[8]/data_i[13] ), .CLK(
        clk), .Q(\read_value_mux[8][13] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[15]  ( .D(\words[8]/data_i[15] ), .CLK(
        clk), .Q(\read_value_mux[8][15] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[17]  ( .D(\words[8]/data_i[17] ), .CLK(
        clk), .Q(\read_value_mux[8][17] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[19]  ( .D(\words[8]/data_i[19] ), .CLK(
        clk), .Q(\read_value_mux[8][19] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[21]  ( .D(\words[8]/data_i[21] ), .CLK(
        clk), .Q(\read_value_mux[8][21] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[23]  ( .D(\words[8]/data_i[23] ), .CLK(
        clk), .Q(\read_value_mux[8][23] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[25]  ( .D(\words[8]/data_i[25] ), .CLK(
        clk), .Q(\read_value_mux[8][25] ) );
  DFFX1_RVT \words[8]/data_ff/data_reg[27]  ( .D(\words[8]/data_i[27] ), .CLK(
        clk), .Q(\read_value_mux[8][27] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[3]  ( .D(\words[11]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[11][3] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[5]  ( .D(\words[11]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[11][5] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[7]  ( .D(\words[11]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[11][7] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[9]  ( .D(\words[11]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[11][9] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[11]  ( .D(\words[11]/data_i[11] ), 
        .CLK(clk), .Q(\read_value_mux[11][11] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[13]  ( .D(\words[11]/data_i[13] ), 
        .CLK(clk), .Q(\read_value_mux[11][13] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[15]  ( .D(\words[11]/data_i[15] ), 
        .CLK(clk), .Q(\read_value_mux[11][15] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[17]  ( .D(\words[11]/data_i[17] ), 
        .CLK(clk), .Q(\read_value_mux[11][17] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[19]  ( .D(\words[11]/data_i[19] ), 
        .CLK(clk), .Q(\read_value_mux[11][19] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[21]  ( .D(\words[11]/data_i[21] ), 
        .CLK(clk), .Q(\read_value_mux[11][21] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[23]  ( .D(\words[11]/data_i[23] ), 
        .CLK(clk), .Q(\read_value_mux[11][23] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[25]  ( .D(\words[11]/data_i[25] ), 
        .CLK(clk), .Q(\read_value_mux[11][25] ) );
  DFFX1_RVT \words[11]/data_ff/data_reg[27]  ( .D(\words[11]/data_i[27] ), 
        .CLK(clk), .Q(\read_value_mux[11][27] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[3]  ( .D(\words[12]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[12][3] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[5]  ( .D(\words[12]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[12][5] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[7]  ( .D(\words[12]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[12][7] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[9]  ( .D(\words[12]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[12][9] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[11]  ( .D(\words[12]/data_i[11] ), 
        .CLK(clk), .Q(\read_value_mux[12][11] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[13]  ( .D(\words[12]/data_i[13] ), 
        .CLK(clk), .Q(\read_value_mux[12][13] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[15]  ( .D(\words[12]/data_i[15] ), 
        .CLK(clk), .Q(\read_value_mux[12][15] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[17]  ( .D(\words[12]/data_i[17] ), 
        .CLK(clk), .Q(\read_value_mux[12][17] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[19]  ( .D(\words[12]/data_i[19] ), 
        .CLK(clk), .Q(\read_value_mux[12][19] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[21]  ( .D(\words[12]/data_i[21] ), 
        .CLK(clk), .Q(\read_value_mux[12][21] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[23]  ( .D(\words[12]/data_i[23] ), 
        .CLK(clk), .Q(\read_value_mux[12][23] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[25]  ( .D(\words[12]/data_i[25] ), 
        .CLK(clk), .Q(\read_value_mux[12][25] ) );
  DFFX1_RVT \words[12]/data_ff/data_reg[27]  ( .D(\words[12]/data_i[27] ), 
        .CLK(clk), .Q(\read_value_mux[12][27] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[3]  ( .D(\words[15]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[15][3] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[5]  ( .D(\words[15]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[15][5] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[7]  ( .D(\words[15]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[15][7] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[9]  ( .D(\words[15]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[15][9] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[11]  ( .D(\words[15]/data_i[11] ), 
        .CLK(clk), .Q(\read_value_mux[15][11] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[13]  ( .D(\words[15]/data_i[13] ), 
        .CLK(clk), .Q(\read_value_mux[15][13] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[15]  ( .D(\words[15]/data_i[15] ), 
        .CLK(clk), .Q(\read_value_mux[15][15] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[17]  ( .D(\words[15]/data_i[17] ), 
        .CLK(clk), .Q(\read_value_mux[15][17] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[19]  ( .D(\words[15]/data_i[19] ), 
        .CLK(clk), .Q(\read_value_mux[15][19] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[21]  ( .D(\words[15]/data_i[21] ), 
        .CLK(clk), .Q(\read_value_mux[15][21] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[23]  ( .D(\words[15]/data_i[23] ), 
        .CLK(clk), .Q(\read_value_mux[15][23] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[25]  ( .D(\words[15]/data_i[25] ), 
        .CLK(clk), .Q(\read_value_mux[15][25] ) );
  DFFX1_RVT \words[15]/data_ff/data_reg[27]  ( .D(\words[15]/data_i[27] ), 
        .CLK(clk), .Q(\read_value_mux[15][27] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[3]  ( .D(\words[16]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[16][3] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[5]  ( .D(\words[16]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[16][5] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[7]  ( .D(\words[16]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[16][7] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[9]  ( .D(\words[16]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[16][9] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[11]  ( .D(\words[16]/data_i[11] ), 
        .CLK(clk), .Q(\read_value_mux[16][11] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[13]  ( .D(\words[16]/data_i[13] ), 
        .CLK(clk), .Q(\read_value_mux[16][13] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[15]  ( .D(\words[16]/data_i[15] ), 
        .CLK(clk), .Q(\read_value_mux[16][15] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[17]  ( .D(\words[16]/data_i[17] ), 
        .CLK(clk), .Q(\read_value_mux[16][17] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[19]  ( .D(\words[16]/data_i[19] ), 
        .CLK(clk), .Q(\read_value_mux[16][19] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[21]  ( .D(\words[16]/data_i[21] ), 
        .CLK(clk), .Q(\read_value_mux[16][21] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[23]  ( .D(\words[16]/data_i[23] ), 
        .CLK(clk), .Q(\read_value_mux[16][23] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[25]  ( .D(\words[16]/data_i[25] ), 
        .CLK(clk), .Q(\read_value_mux[16][25] ) );
  DFFX1_RVT \words[16]/data_ff/data_reg[27]  ( .D(\words[16]/data_i[27] ), 
        .CLK(clk), .Q(\read_value_mux[16][27] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[3]  ( .D(\words[20]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[20][3] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[5]  ( .D(\words[20]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[20][5] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[7]  ( .D(\words[20]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[20][7] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[9]  ( .D(\words[20]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[20][9] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[11]  ( .D(\words[20]/data_i[11] ), 
        .CLK(clk), .Q(\read_value_mux[20][11] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[13]  ( .D(\words[20]/data_i[13] ), 
        .CLK(clk), .Q(\read_value_mux[20][13] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[15]  ( .D(\words[20]/data_i[15] ), 
        .CLK(clk), .Q(\read_value_mux[20][15] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[17]  ( .D(\words[20]/data_i[17] ), 
        .CLK(clk), .Q(\read_value_mux[20][17] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[19]  ( .D(\words[20]/data_i[19] ), 
        .CLK(clk), .Q(\read_value_mux[20][19] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[21]  ( .D(\words[20]/data_i[21] ), 
        .CLK(clk), .Q(\read_value_mux[20][21] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[23]  ( .D(\words[20]/data_i[23] ), 
        .CLK(clk), .Q(\read_value_mux[20][23] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[25]  ( .D(\words[20]/data_i[25] ), 
        .CLK(clk), .Q(\read_value_mux[20][25] ) );
  DFFX1_RVT \words[20]/data_ff/data_reg[27]  ( .D(\words[20]/data_i[27] ), 
        .CLK(clk), .Q(\read_value_mux[20][27] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[3]  ( .D(\words[23]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[23][3] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[5]  ( .D(\words[23]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[23][5] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[7]  ( .D(\words[23]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[23][7] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[9]  ( .D(\words[23]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[23][9] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[11]  ( .D(\words[23]/data_i[11] ), 
        .CLK(clk), .Q(\read_value_mux[23][11] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[13]  ( .D(\words[23]/data_i[13] ), 
        .CLK(clk), .Q(\read_value_mux[23][13] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[15]  ( .D(\words[23]/data_i[15] ), 
        .CLK(clk), .Q(\read_value_mux[23][15] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[17]  ( .D(\words[23]/data_i[17] ), 
        .CLK(clk), .Q(\read_value_mux[23][17] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[19]  ( .D(\words[23]/data_i[19] ), 
        .CLK(clk), .Q(\read_value_mux[23][19] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[21]  ( .D(\words[23]/data_i[21] ), 
        .CLK(clk), .Q(\read_value_mux[23][21] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[23]  ( .D(\words[23]/data_i[23] ), 
        .CLK(clk), .Q(\read_value_mux[23][23] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[25]  ( .D(\words[23]/data_i[25] ), 
        .CLK(clk), .Q(\read_value_mux[23][25] ) );
  DFFX1_RVT \words[23]/data_ff/data_reg[27]  ( .D(\words[23]/data_i[27] ), 
        .CLK(clk), .Q(\read_value_mux[23][27] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[3]  ( .D(\words[24]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[24][3] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[5]  ( .D(\words[24]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[24][5] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[7]  ( .D(\words[24]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[24][7] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[9]  ( .D(\words[24]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[24][9] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[11]  ( .D(\words[24]/data_i[11] ), 
        .CLK(clk), .Q(\read_value_mux[24][11] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[13]  ( .D(\words[24]/data_i[13] ), 
        .CLK(clk), .Q(\read_value_mux[24][13] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[15]  ( .D(\words[24]/data_i[15] ), 
        .CLK(clk), .Q(\read_value_mux[24][15] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[17]  ( .D(\words[24]/data_i[17] ), 
        .CLK(clk), .Q(\read_value_mux[24][17] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[19]  ( .D(\words[24]/data_i[19] ), 
        .CLK(clk), .Q(\read_value_mux[24][19] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[21]  ( .D(\words[24]/data_i[21] ), 
        .CLK(clk), .Q(\read_value_mux[24][21] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[23]  ( .D(\words[24]/data_i[23] ), 
        .CLK(clk), .Q(\read_value_mux[24][23] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[25]  ( .D(\words[24]/data_i[25] ), 
        .CLK(clk), .Q(\read_value_mux[24][25] ) );
  DFFX1_RVT \words[24]/data_ff/data_reg[27]  ( .D(\words[24]/data_i[27] ), 
        .CLK(clk), .Q(\read_value_mux[24][27] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[3]  ( .D(\words[27]/data_i[3] ), .CLK(
        clk), .Q(\read_value_mux[27][3] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[5]  ( .D(\words[27]/data_i[5] ), .CLK(
        clk), .Q(\read_value_mux[27][5] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[7]  ( .D(\words[27]/data_i[7] ), .CLK(
        clk), .Q(\read_value_mux[27][7] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[9]  ( .D(\words[27]/data_i[9] ), .CLK(
        clk), .Q(\read_value_mux[27][9] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[11]  ( .D(\words[27]/data_i[11] ), 
        .CLK(clk), .Q(\read_value_mux[27][11] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[13]  ( .D(\words[27]/data_i[13] ), 
        .CLK(clk), .Q(\read_value_mux[27][13] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[15]  ( .D(\words[27]/data_i[15] ), 
        .CLK(clk), .Q(\read_value_mux[27][15] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[17]  ( .D(\words[27]/data_i[17] ), 
        .CLK(clk), .Q(\read_value_mux[27][17] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[19]  ( .D(\words[27]/data_i[19] ), 
        .CLK(clk), .Q(\read_value_mux[27][19] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[21]  ( .D(\words[27]/data_i[21] ), 
        .CLK(clk), .Q(\read_value_mux[27][21] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[23]  ( .D(\words[27]/data_i[23] ), 
        .CLK(clk), .Q(\read_value_mux[27][23] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[25]  ( .D(\words[27]/data_i[25] ), 
        .CLK(clk), .Q(\read_value_mux[27][25] ) );
  DFFX1_RVT \words[27]/data_ff/data_reg[27]  ( .D(\words[27]/data_i[27] ), 
        .CLK(clk), .Q(\read_value_mux[27][27] ) );
  AO221X1_RVT U2478 ( .A1(1'b1), .A2(read_index[2]), .A3(n1777), .A4(
        \words[0]/valid_o ), .A5(n1774), .Y(n1501) );
  AO221X1_RVT U2479 ( .A1(1'b1), .A2(n3107), .A3(n3106), .A4(n1492), .A5(n3105), .Y(n1494) );
  AO221X1_RVT U2480 ( .A1(1'b1), .A2(n3004), .A3(n3012), .A4(n1481), .A5(n3006), .Y(n2988) );
  OA221X1_RVT U2481 ( .A1(1'b0), .A2(n3011), .A3(n2991), .A4(n2990), .A5(n3009), .Y(n2987) );
  INVX1_RVT U2482 ( .A(search_data[17]), .Y(n1715) );
  INVX1_RVT U2483 ( .A(search_data[9]), .Y(n1737) );
  INVX1_RVT U2484 ( .A(reset), .Y(n3085) );
  NAND4X0_RVT U2486 ( .A1(n2985), .A2(n2984), .A3(n2996), .A4(n2986), .Y(n1480) );
  OAI21X1_RVT U2487 ( .A1(n3008), .A2(n2987), .A3(n1480), .Y(n1481) );
  NOR4X0_RVT U2489 ( .A1(n3007), .A2(n3006), .A3(n2976), .A4(n2953), .Y(n1483)
         );
  AO221X1_RVT U2490 ( .A1(n3100), .A2(n2907), .A3(n3100), .A4(n2980), .A5(
        n2961), .Y(n1484) );
  AO21X1_RVT U2491 ( .A1(n2954), .A2(n1484), .A3(n2955), .Y(n1485) );
  INVX0_RVT U2492 ( .A(n3006), .Y(n1486) );
  OA221X1_RVT U2493 ( .A1(n3008), .A2(n2978), .A3(n3008), .A4(n3011), .A5(
        n3012), .Y(n1487) );
  AO221X1_RVT U2494 ( .A1(n1486), .A2(n3004), .A3(n1486), .A4(n1487), .A5(
        n3005), .Y(n1488) );
  AO22X1_RVT U2495 ( .A1(n1483), .A2(n1485), .A3(n2989), .A4(n1488), .Y(
        search_index[0]) );
  AO21X1_RVT U2496 ( .A1(n1689), .A2(n1690), .A3(n2988), .Y(n1489) );
  INVX0_RVT U2497 ( .A(n3005), .Y(n1490) );
  AND3X1_RVT U2498 ( .A1(n2989), .A2(n1489), .A3(n1490), .Y(search_index[1])
         );
  NAND4X0_RVT U2499 ( .A1(n3098), .A2(n3099), .A3(n3100), .A4(n3101), .Y(n1491) );
  NAND4X0_RVT U2500 ( .A1(n3102), .A2(n3103), .A3(n3104), .A4(n1491), .Y(n1492) );
  OA221X1_RVT U2502 ( .A1(n3110), .A2(n3109), .A3(n3110), .A4(n1494), .A5(
        n3108), .Y(search_index[2]) );
  AO21X1_RVT U2503 ( .A1(\words[8]/valid_o ), .A2(n1777), .A3(n1688), .Y(n1495) );
  NAND2X0_RVT U2504 ( .A1(n1778), .A2(\words[14]/valid_o ), .Y(n1496) );
  NAND4X0_RVT U2505 ( .A1(read_index[2]), .A2(n1772), .A3(n1773), .A4(n1496), 
        .Y(n1497) );
  OA221X1_RVT U2506 ( .A1(n1495), .A2(n1778), .A3(n1495), .A4(
        \words[10]/valid_o ), .A5(n1497), .Y(n1498) );
  INVX0_RVT U2507 ( .A(read_index[3]), .Y(n1499) );
  INVX0_RVT U2509 ( .A(read_index[2]), .Y(n1502) );
  AO22X1_RVT U2510 ( .A1(n1776), .A2(\words[5]/valid_o ), .A3(n1775), .A4(
        \words[7]/valid_o ), .Y(n1503) );
  AO22X1_RVT U2511 ( .A1(n1777), .A2(\words[4]/valid_o ), .A3(n1778), .A4(
        \words[6]/valid_o ), .Y(n1504) );
  OR3X1_RVT U2512 ( .A1(n1502), .A2(n1503), .A3(n1504), .Y(n1505) );
  OA221X1_RVT U2513 ( .A1(n1501), .A2(n1778), .A3(n1501), .A4(
        \words[2]/valid_o ), .A5(n1505), .Y(n1506) );
  AO22X1_RVT U2514 ( .A1(read_index[3]), .A2(n1498), .A3(n1499), .A4(n1506), 
        .Y(n1507) );
  INVX0_RVT U2515 ( .A(read_index[4]), .Y(n1508) );
  OA22X1_RVT U2516 ( .A1(n1779), .A2(\words[31]/valid_o ), .A3(n1780), .A4(
        \words[29]/valid_o ), .Y(n1509) );
  OA22X1_RVT U2517 ( .A1(n1782), .A2(\words[28]/valid_o ), .A3(n1781), .A4(
        \words[30]/valid_o ), .Y(n1510) );
  NAND3X0_RVT U2518 ( .A1(read_index[2]), .A2(n1509), .A3(n1510), .Y(n1511) );
  OA22X1_RVT U2519 ( .A1(n1779), .A2(\words[27]/valid_o ), .A3(n1780), .A4(
        \words[25]/valid_o ), .Y(n1512) );
  OA22X1_RVT U2520 ( .A1(n1782), .A2(\words[24]/valid_o ), .A3(n1781), .A4(
        \words[26]/valid_o ), .Y(n1513) );
  NAND3X0_RVT U2521 ( .A1(n1512), .A2(n1513), .A3(n1502), .Y(n1514) );
  NAND2X0_RVT U2522 ( .A1(n1511), .A2(n1514), .Y(n1515) );
  OA22X1_RVT U2523 ( .A1(n1779), .A2(\words[23]/valid_o ), .A3(n1780), .A4(
        \words[21]/valid_o ), .Y(n1516) );
  OA22X1_RVT U2524 ( .A1(n1782), .A2(\words[20]/valid_o ), .A3(n1781), .A4(
        \words[22]/valid_o ), .Y(n1517) );
  NAND3X0_RVT U2525 ( .A1(read_index[2]), .A2(n1516), .A3(n1517), .Y(n1518) );
  OA22X1_RVT U2526 ( .A1(n1779), .A2(\words[19]/valid_o ), .A3(n1780), .A4(
        \words[17]/valid_o ), .Y(n1519) );
  OA22X1_RVT U2527 ( .A1(n1782), .A2(\words[16]/valid_o ), .A3(n1781), .A4(
        \words[18]/valid_o ), .Y(n1520) );
  NAND3X0_RVT U2528 ( .A1(n1519), .A2(n1520), .A3(n1502), .Y(n1521) );
  NAND2X0_RVT U2529 ( .A1(n1518), .A2(n1521), .Y(n1522) );
  AO22X1_RVT U2530 ( .A1(read_index[3]), .A2(n1515), .A3(n1499), .A4(n1522), 
        .Y(n1523) );
  OA221X1_RVT U2531 ( .A1(read_index[4]), .A2(n1507), .A3(n1508), .A4(n1523), 
        .A5(read), .Y(read_valid) );
  NBUFFX8_RVT U2532 ( .A(n2940), .Y(n1738) );
  IBUFFX8_RVT U2533 ( .A(search_data[6]), .Y(n2940) );
  NBUFFX4_RVT U2534 ( .A(n1741), .Y(n1740) );
  NBUFFX4_RVT U2535 ( .A(n1741), .Y(n1739) );
  IBUFFX8_RVT U2536 ( .A(search_data[7]), .Y(n1741) );
  IBUFFX16_RVT U2537 ( .A(search_data[3]), .Y(n1750) );
  INVX0_RVT U2538 ( .A(n3014), .Y(n3115) );
  INVX0_RVT U2539 ( .A(n3015), .Y(n3111) );
  INVX0_RVT U2540 ( .A(n3110), .Y(n3013) );
  INVX0_RVT U2541 ( .A(n3098), .Y(n3003) );
  INVX0_RVT U2542 ( .A(n3107), .Y(n2995) );
  INVX0_RVT U2543 ( .A(n2958), .Y(n2431) );
  AND2X1_RVT U2544 ( .A1(n3074), .A2(n3087), .Y(n3075) );
  AND2X1_RVT U2545 ( .A1(n3074), .A2(n3095), .Y(n3044) );
  AND2X1_RVT U2546 ( .A1(n3074), .A2(n3080), .Y(n3065) );
  AND2X1_RVT U2547 ( .A1(n3091), .A2(n3074), .Y(n3019) );
  AND2X1_RVT U2548 ( .A1(n3080), .A2(n3041), .Y(n3038) );
  NOR3X1_RVT U2549 ( .A1(write_index[2]), .A2(write_index[3]), .A3(n3018), .Y(
        n3074) );
  AND2X1_RVT U2550 ( .A1(n3096), .A2(n3095), .Y(n3097) );
  AND2X1_RVT U2551 ( .A1(n3080), .A2(n3032), .Y(n3029) );
  AND2X1_RVT U2552 ( .A1(n3087), .A2(n3032), .Y(n3033) );
  AND2X1_RVT U2553 ( .A1(n3095), .A2(n3041), .Y(n3037) );
  AND2X1_RVT U2554 ( .A1(n3091), .A2(n3096), .Y(n3092) );
  AND2X1_RVT U2555 ( .A1(n3032), .A2(n3095), .Y(n3028) );
  AND2X1_RVT U2556 ( .A1(n3091), .A2(n3052), .Y(n3046) );
  AND2X1_RVT U2557 ( .A1(n3080), .A2(n3052), .Y(n3049) );
  AND2X1_RVT U2558 ( .A1(n3096), .A2(n3080), .Y(n3021) );
  AND2X1_RVT U2559 ( .A1(n3087), .A2(n3052), .Y(n3053) );
  AND2X1_RVT U2560 ( .A1(n3096), .A2(n3087), .Y(n3023) );
  AND2X1_RVT U2561 ( .A1(n3095), .A2(n3052), .Y(n3048) );
  AND2X1_RVT U2562 ( .A1(n3091), .A2(n3032), .Y(n3024) );
  AO21X1_RVT U2563 ( .A1(n3088), .A2(n3086), .A3(reset), .Y(n3083) );
  AO21X1_RVT U2564 ( .A1(n3060), .A2(n3069), .A3(reset), .Y(n3059) );
  AO21X1_RVT U2565 ( .A1(n3088), .A2(n3070), .A3(reset), .Y(n3031) );
  AO21X1_RVT U2566 ( .A1(n3088), .A2(n3035), .A3(reset), .Y(n3073) );
  AND2X1_RVT U2567 ( .A1(n3091), .A2(n3041), .Y(n3036) );
  AO21X1_RVT U2568 ( .A1(n3088), .A2(n3060), .A3(reset), .Y(n3094) );
  AO21X1_RVT U2569 ( .A1(n3069), .A2(n3086), .A3(reset), .Y(n3051) );
  AND2X1_RVT U2570 ( .A1(n3087), .A2(n3041), .Y(n3042) );
  AO21X1_RVT U2571 ( .A1(n3070), .A2(n3069), .A3(reset), .Y(n3068) );
  OR2X1_RVT U2572 ( .A1(n3026), .A2(write_index[1]), .Y(n3027) );
  OR2X1_RVT U2573 ( .A1(write_index[1]), .A2(write_index[0]), .Y(n3017) );
  INVX0_RVT U2574 ( .A(read_index[0]), .Y(n1771) );
  NOR2X1_RVT U2575 ( .A1(write_index[2]), .A2(write_index[3]), .Y(n3035) );
  INVX0_RVT U2576 ( .A(read_index[1]), .Y(n1769) );
  NBUFFX8_RVT U2577 ( .A(n1749), .Y(n1524) );
  NBUFFX8_RVT U2578 ( .A(n1747), .Y(n1525) );
  NBUFFX4_RVT U2579 ( .A(n2942), .Y(n1526) );
  NBUFFX4_RVT U2580 ( .A(n2934), .Y(n1527) );
  NBUFFX4_RVT U2581 ( .A(n1731), .Y(n1528) );
  NBUFFX4_RVT U2582 ( .A(n1729), .Y(n1529) );
  NBUFFX8_RVT U2583 ( .A(n1726), .Y(n1530) );
  NBUFFX4_RVT U2584 ( .A(n2931), .Y(n1531) );
  NBUFFX4_RVT U2585 ( .A(n2929), .Y(n1532) );
  NBUFFX4_RVT U2586 ( .A(n2923), .Y(n1533) );
  NBUFFX4_RVT U2587 ( .A(n1709), .Y(n1534) );
  NBUFFX4_RVT U2588 ( .A(n1707), .Y(n1535) );
  NBUFFX4_RVT U2589 ( .A(n1704), .Y(n1536) );
  NBUFFX4_RVT U2590 ( .A(n2920), .Y(n1537) );
  NBUFFX8_RVT U2591 ( .A(n1700), .Y(n1538) );
  NBUFFX4_RVT U2592 ( .A(n2918), .Y(n1539) );
  NBUFFX8_RVT U2593 ( .A(n1697), .Y(n1540) );
  NBUFFX4_RVT U2594 ( .A(n2912), .Y(n1541) );
  NBUFFX8_RVT U2595 ( .A(n1694), .Y(n1542) );
  NBUFFX4_RVT U2596 ( .A(n1693), .Y(n1543) );
  NAND2X0_RVT U2597 ( .A1(n3090), .A2(n3059), .Y(n1677) );
  NAND2X0_RVT U2598 ( .A1(n3090), .A2(n3083), .Y(n1679) );
  NAND2X0_RVT U2599 ( .A1(n3090), .A2(n3068), .Y(n1678) );
  NAND2X0_RVT U2600 ( .A1(n3017), .A2(n3085), .Y(n3090) );
  NAND2X0_RVT U2601 ( .A1(n3079), .A2(n3083), .Y(n3082) );
  NAND2X0_RVT U2602 ( .A1(n3084), .A2(n3083), .Y(n1634) );
  NAND2X0_RVT U2603 ( .A1(n3084), .A2(n3068), .Y(n3072) );
  NAND2X0_RVT U2604 ( .A1(n3079), .A2(n3068), .Y(n3067) );
  NAND2X0_RVT U2605 ( .A1(n3084), .A2(n3059), .Y(n1633) );
  NAND2X0_RVT U2606 ( .A1(n3079), .A2(n3059), .Y(n3058) );
  NAND2X0_RVT U2607 ( .A1(n3093), .A2(n3068), .Y(n3064) );
  NAND2X0_RVT U2608 ( .A1(n3093), .A2(n3059), .Y(n1683) );
  NAND2X0_RVT U2609 ( .A1(n3093), .A2(n3083), .Y(n1684) );
  NAND2X0_RVT U2610 ( .A1(n3085), .A2(n3022), .Y(n3084) );
  NAND2X0_RVT U2611 ( .A1(n3085), .A2(n3020), .Y(n3079) );
  NAND2X0_RVT U2612 ( .A1(n3085), .A2(n3027), .Y(n3093) );
  AND2X1_RVT U2613 ( .A1(write), .A2(n3016), .Y(n3088) );
  OA221X1_RVT U2614 ( .A1(n3014), .A2(n3112), .A3(n3014), .A4(n3015), .A5(
        n3114), .Y(search_index[3]) );
  NAND2X0_RVT U2615 ( .A1(n3090), .A2(n3094), .Y(n1680) );
  NAND2X0_RVT U2616 ( .A1(n3090), .A2(n3031), .Y(n3025) );
  NAND2X0_RVT U2617 ( .A1(n3090), .A2(n3073), .Y(n1675) );
  NAND2X0_RVT U2618 ( .A1(n3090), .A2(n3051), .Y(n3047) );
  NAND2X0_RVT U2619 ( .A1(n3090), .A2(n3040), .Y(n1676) );
  NAND2X0_RVT U2620 ( .A1(n3079), .A2(n3051), .Y(n3050) );
  NAND2X0_RVT U2621 ( .A1(n3084), .A2(n3031), .Y(n1631) );
  NAND2X0_RVT U2622 ( .A1(n3079), .A2(n3031), .Y(n3030) );
  NAND2X0_RVT U2623 ( .A1(n3084), .A2(n3051), .Y(n3054) );
  NAND2X0_RVT U2624 ( .A1(n3084), .A2(n3040), .Y(n3043) );
  NAND2X0_RVT U2625 ( .A1(n3079), .A2(n3040), .Y(n3039) );
  NAND2X0_RVT U2626 ( .A1(n3093), .A2(n3051), .Y(n1682) );
  NAND2X0_RVT U2627 ( .A1(n3093), .A2(n3040), .Y(n1681) );
  NAND2X0_RVT U2628 ( .A1(n3094), .A2(n3084), .Y(n1686) );
  NAND2X0_RVT U2629 ( .A1(n3073), .A2(n3084), .Y(n3076) );
  NAND2X0_RVT U2630 ( .A1(n3094), .A2(n3079), .Y(n1685) );
  NAND2X0_RVT U2631 ( .A1(n3073), .A2(n3079), .Y(n1687) );
  NAND2X0_RVT U2632 ( .A1(n3094), .A2(n3093), .Y(n1635) );
  NAND2X0_RVT U2633 ( .A1(n3073), .A2(n3093), .Y(n1632) );
  NAND2X0_RVT U2634 ( .A1(n3031), .A2(n3093), .Y(n1630) );
  NOR2X0_RVT U2635 ( .A1(n3045), .A2(write_index[3]), .Y(n3086) );
  AND2X1_RVT U2636 ( .A1(write_index[3]), .A2(n3045), .Y(n3060) );
  INVX1_RVT U2637 ( .A(n3027), .Y(n3095) );
  INVX1_RVT U2638 ( .A(search_data[25]), .Y(n1697) );
  AND4X1_RVT U2639 ( .A1(n3091), .A2(n3060), .A3(n3069), .A4(n3085), .Y(n3055)
         );
  AND4X1_RVT U2640 ( .A1(n3091), .A2(n3088), .A3(n3086), .A4(n3085), .Y(n3077)
         );
  AND4X1_RVT U2641 ( .A1(n3091), .A2(n3070), .A3(n3069), .A4(n3085), .Y(n3062)
         );
  INVX1_RVT U2642 ( .A(n3017), .Y(n3091) );
  AND4X1_RVT U2643 ( .A1(n3088), .A2(n3080), .A3(n3086), .A4(n3085), .Y(n3081)
         );
  AND4X1_RVT U2644 ( .A1(n3088), .A2(n3087), .A3(n3086), .A4(n3085), .Y(n3089)
         );
  AND4X1_RVT U2645 ( .A1(n3087), .A2(n3070), .A3(n3069), .A4(n3085), .Y(n3071)
         );
  AND4X1_RVT U2646 ( .A1(n3080), .A2(n3070), .A3(n3069), .A4(n3085), .Y(n3066)
         );
  AND4X1_RVT U2647 ( .A1(n3060), .A2(n3087), .A3(n3069), .A4(n3085), .Y(n3061)
         );
  AND4X1_RVT U2648 ( .A1(n3060), .A2(n3080), .A3(n3069), .A4(n3085), .Y(n3057)
         );
  AND4X1_RVT U2649 ( .A1(n3070), .A2(n3095), .A3(n3069), .A4(n3085), .Y(n3063)
         );
  AND4X1_RVT U2650 ( .A1(n3060), .A2(n3095), .A3(n3069), .A4(n3085), .Y(n3056)
         );
  AND4X1_RVT U2651 ( .A1(n3088), .A2(n3095), .A3(n3086), .A4(n3085), .Y(n3078)
         );
  INVX1_RVT U2652 ( .A(n3020), .Y(n3080) );
  OR4X1_RVT U2653 ( .A1(n2142), .A2(n2141), .A3(n2140), .A4(n2139), .Y(n2994)
         );
  INVX1_RVT U2654 ( .A(search_data[13]), .Y(n1726) );
  INVX1_RVT U2655 ( .A(search_data[23]), .Y(n1700) );
  INVX1_RVT U2656 ( .A(search_data[27]), .Y(n1694) );
  NAND2X0_RVT U2657 ( .A1(n3085), .A2(n3034), .Y(n3040) );
  AND2X1_RVT U2658 ( .A1(write_index[4]), .A2(write), .Y(n3069) );
  AND3X1_RVT U2659 ( .A1(n3115), .A2(n3114), .A3(n3113), .Y(search_index[4])
         );
  INVX1_RVT U2660 ( .A(search_data[30]), .Y(n1764) );
  INVX1_RVT U2661 ( .A(search_data[28]), .Y(n1758) );
  OR4X1_RVT U2662 ( .A1(n2034), .A2(n2033), .A3(n2032), .A4(n2031), .Y(n3012)
         );
  NAND2X0_RVT U2663 ( .A1(write_index[1]), .A2(n3026), .Y(n3020) );
  INVX1_RVT U2664 ( .A(write_index[2]), .Y(n3045) );
  AND2X1_RVT U2665 ( .A1(write_index[2]), .A2(write_index[3]), .Y(n3070) );
  OR4X1_RVT U2666 ( .A1(n2690), .A2(n2689), .A3(n2688), .A4(n2687), .Y(n3100)
         );
  OR4X1_RVT U2667 ( .A1(n1998), .A2(n1997), .A3(n1996), .A4(n1995), .Y(n3011)
         );
  INVX1_RVT U2668 ( .A(search_data[2]), .Y(n1749) );
  INVX1_RVT U2669 ( .A(search_data[4]), .Y(n2942) );
  INVX1_RVT U2670 ( .A(search_data[5]), .Y(n1747) );
  INVX1_RVT U2671 ( .A(search_data[8]), .Y(n2934) );
  INVX1_RVT U2672 ( .A(search_data[10]), .Y(n1729) );
  INVX1_RVT U2673 ( .A(search_data[11]), .Y(n1731) );
  INVX1_RVT U2674 ( .A(search_data[12]), .Y(n2931) );
  INVX1_RVT U2675 ( .A(search_data[14]), .Y(n2929) );
  INVX1_RVT U2676 ( .A(search_data[15]), .Y(n1723) );
  INVX1_RVT U2677 ( .A(search_data[16]), .Y(n2923) );
  INVX1_RVT U2678 ( .A(search_data[18]), .Y(n1707) );
  INVX1_RVT U2679 ( .A(search_data[19]), .Y(n1709) );
  INVX1_RVT U2680 ( .A(search_data[20]), .Y(n2920) );
  INVX1_RVT U2681 ( .A(search_data[21]), .Y(n1704) );
  INVX1_RVT U2682 ( .A(search_data[22]), .Y(n2918) );
  INVX1_RVT U2683 ( .A(search_data[24]), .Y(n2912) );
  INVX1_RVT U2684 ( .A(search_data[26]), .Y(n1693) );
  INVX1_RVT U2685 ( .A(search_data[30]), .Y(n1763) );
  INVX1_RVT U2686 ( .A(search_data[28]), .Y(n1757) );
  INVX1_RVT U2687 ( .A(write_index[0]), .Y(n3026) );
  INVX1_RVT U2688 ( .A(write_index[4]), .Y(n3016) );
  NOR2X0_RVT U2689 ( .A1(n2958), .A2(n2957), .Y(n3104) );
  OR4X1_RVT U2690 ( .A1(n2540), .A2(n2539), .A3(n2538), .A4(n2537), .Y(n2971)
         );
  INVX1_RVT U2691 ( .A(search_data[31]), .Y(n1767) );
  INVX1_RVT U2692 ( .A(search_data[29]), .Y(n1761) );
  OR4X1_RVT U2693 ( .A1(n2106), .A2(n2105), .A3(n2104), .A4(n2103), .Y(n2975)
         );
  INVX1_RVT U2694 ( .A(search_data[0]), .Y(n1752) );
  INVX1_RVT U2695 ( .A(search_data[1]), .Y(n1755) );
  INVX1_RVT U2696 ( .A(search_data[31]), .Y(n1768) );
  INVX1_RVT U2697 ( .A(search_data[29]), .Y(n1762) );
  INVX1_RVT U2698 ( .A(search_data[31]), .Y(n1766) );
  INVX1_RVT U2699 ( .A(search_data[29]), .Y(n1760) );
  INVX1_RVT U2700 ( .A(n3022), .Y(n3087) );
  NAND4X0_RVT U2701 ( .A1(n3114), .A2(n3115), .A3(n3112), .A4(n3111), .Y(
        search_valid) );
  AND2X1_RVT U2702 ( .A1(n2963), .A2(n2962), .Y(n3101) );
  OR2X1_RVT U2703 ( .A1(n2977), .A2(n2976), .Y(n2990) );
  OR4X1_RVT U2704 ( .A1(n2214), .A2(n2213), .A3(n2212), .A4(n2211), .Y(n2985)
         );
  INVX1_RVT U2705 ( .A(search_data[1]), .Y(n1756) );
  INVX1_RVT U2706 ( .A(search_data[1]), .Y(n1754) );
  AND2X1_RVT U2707 ( .A1(n3108), .A2(n3013), .Y(n3114) );
  OR4X1_RVT U2708 ( .A1(n2870), .A2(n2869), .A3(n2868), .A4(n2867), .Y(n3002)
         );
  OR4X1_RVT U2709 ( .A1(n2651), .A2(n2650), .A3(n2649), .A4(n2648), .Y(n2962)
         );
  INVX1_RVT U2710 ( .A(n2654), .Y(n3103) );
  NBUFFX2_RVT U2711 ( .A(n1731), .Y(n1730) );
  NBUFFX2_RVT U2712 ( .A(n1709), .Y(n1708) );
  NBUFFX2_RVT U2713 ( .A(n1704), .Y(n1703) );
  AND4X1_RVT U2714 ( .A1(write_index[4]), .A2(write), .A3(n3086), .A4(n3085), 
        .Y(n3052) );
  AND4X1_RVT U2715 ( .A1(write_index[4]), .A2(write), .A3(n3035), .A4(n3085), 
        .Y(n3041) );
  NAND2X0_RVT U2716 ( .A1(write_index[1]), .A2(write_index[0]), .Y(n3022) );
  AND4X1_RVT U2717 ( .A1(n3088), .A2(write_index[3]), .A3(n3085), .A4(n3045), 
        .Y(n3096) );
  NAND2X0_RVT U2718 ( .A1(n3088), .A2(n3085), .Y(n3018) );
  AND4X1_RVT U2719 ( .A1(n3088), .A2(write_index[2]), .A3(write_index[3]), 
        .A4(n3085), .Y(n3032) );
  AND4X1_RVT U2720 ( .A1(n3104), .A2(n3106), .A3(n3103), .A4(n3102), .Y(n3112)
         );
  INVX1_RVT U2721 ( .A(n1781), .Y(n1778) );
  OR2X1_RVT U2722 ( .A1(read_index[2]), .A2(n1770), .Y(n1688) );
  INVX1_RVT U2723 ( .A(n1779), .Y(n1775) );
  INVX1_RVT U2724 ( .A(n1780), .Y(n1776) );
  INVX1_RVT U2725 ( .A(n1782), .Y(n1777) );
  OR2X1_RVT U2726 ( .A1(n3107), .A2(n2972), .Y(n1690) );
  NOR4X1_RVT U2727 ( .A1(n2977), .A2(n2976), .A3(n3008), .A4(n3105), .Y(n2986)
         );
  INVX1_RVT U2728 ( .A(n2980), .Y(n3099) );
  INVX1_RVT U2729 ( .A(n2965), .Y(n3000) );
  INVX1_RVT U2730 ( .A(n2964), .Y(n3001) );
  INVX1_RVT U2731 ( .A(n2961), .Y(n2963) );
  INVX1_RVT U2732 ( .A(n2960), .Y(n3102) );
  INVX1_RVT U2733 ( .A(n2959), .Y(n2996) );
  INVX1_RVT U2734 ( .A(n2979), .Y(n2997) );
  INVX1_RVT U2735 ( .A(n2956), .Y(n2993) );
  INVX1_RVT U2736 ( .A(n2973), .Y(n2974) );
  INVX1_RVT U2737 ( .A(n2990), .Y(n2992) );
  INVX1_RVT U2738 ( .A(n2969), .Y(n2970) );
  INVX1_RVT U2739 ( .A(n2978), .Y(n3009) );
  INVX1_RVT U2740 ( .A(n3008), .Y(n3010) );
  NOR4X1_RVT U2741 ( .A1(n3007), .A2(n3006), .A3(n3005), .A4(n3004), .Y(n3108)
         );
  NOR4X1_RVT U2742 ( .A1(n2952), .A2(n2951), .A3(n2950), .A4(n2949), .Y(n2976)
         );
  NOR4X1_RVT U2743 ( .A1(n2906), .A2(n2905), .A3(n2904), .A4(n2903), .Y(n2961)
         );
  NOR4X1_RVT U2744 ( .A1(n2798), .A2(n2797), .A3(n2796), .A4(n2795), .Y(n2965)
         );
  NOR4X1_RVT U2745 ( .A1(n2762), .A2(n2761), .A3(n2760), .A4(n2759), .Y(n2964)
         );
  NOR4X1_RVT U2746 ( .A1(n2726), .A2(n2725), .A3(n2724), .A4(n2723), .Y(n2980)
         );
  NOR4X1_RVT U2747 ( .A1(n2654), .A2(n2958), .A3(n2653), .A4(n2652), .Y(n2954)
         );
  NOR4X1_RVT U2748 ( .A1(n2614), .A2(n2613), .A3(n2612), .A4(n2611), .Y(n2977)
         );
  NOR4X1_RVT U2749 ( .A1(n2577), .A2(n2576), .A3(n2575), .A4(n2574), .Y(n2973)
         );
  NOR4X1_RVT U2750 ( .A1(n2504), .A2(n2503), .A3(n2502), .A4(n2501), .Y(n2959)
         );
  NOR4X1_RVT U2751 ( .A1(n2467), .A2(n2466), .A3(n2465), .A4(n2464), .Y(n2969)
         );
  NBUFFX2_RVT U2752 ( .A(n1723), .Y(n1720) );
  NOR4X1_RVT U2753 ( .A1(n2430), .A2(n2429), .A3(n2428), .A4(n2427), .Y(n2958)
         );
  NOR4X1_RVT U2754 ( .A1(n2394), .A2(n2393), .A3(n2392), .A4(n2391), .Y(n2654)
         );
  NOR4X1_RVT U2755 ( .A1(n2358), .A2(n2357), .A3(n2356), .A4(n2355), .Y(n2960)
         );
  NOR4X1_RVT U2756 ( .A1(n2322), .A2(n2321), .A3(n2320), .A4(n2319), .Y(n2957)
         );
  NOR4X1_RVT U2757 ( .A1(n2286), .A2(n2285), .A3(n2284), .A4(n2283), .Y(n2979)
         );
  INVX1_RVT U2758 ( .A(n2653), .Y(n2998) );
  NOR4X1_RVT U2759 ( .A1(n2178), .A2(n2177), .A3(n2176), .A4(n2175), .Y(n2956)
         );
  NBUFFX2_RVT U2760 ( .A(n1747), .Y(n1745) );
  NBUFFX2_RVT U2761 ( .A(n1723), .Y(n1721) );
  NOR4X1_RVT U2762 ( .A1(n2070), .A2(n2069), .A3(n2068), .A4(n2067), .Y(n3005)
         );
  NOR4X1_RVT U2763 ( .A1(n1962), .A2(n1961), .A3(n1960), .A4(n1959), .Y(n2978)
         );
  NOR4X1_RVT U2764 ( .A1(n1926), .A2(n1925), .A3(n1924), .A4(n1923), .Y(n3008)
         );
  NBUFFX2_RVT U2765 ( .A(n1729), .Y(n1728) );
  NBUFFX2_RVT U2766 ( .A(n2923), .Y(n1711) );
  NBUFFX2_RVT U2767 ( .A(n1707), .Y(n1706) );
  NBUFFX2_RVT U2768 ( .A(n2920), .Y(n1702) );
  NBUFFX2_RVT U2769 ( .A(n1693), .Y(n1692) );
  NOR4X1_RVT U2770 ( .A1(n1890), .A2(n1889), .A3(n1888), .A4(n1887), .Y(n3004)
         );
  NBUFFX2_RVT U2771 ( .A(n1749), .Y(n1748) );
  NBUFFX2_RVT U2772 ( .A(n2942), .Y(n1743) );
  NBUFFX2_RVT U2773 ( .A(n2934), .Y(n1733) );
  NBUFFX2_RVT U2774 ( .A(n2931), .Y(n1725) );
  NBUFFX2_RVT U2775 ( .A(n2929), .Y(n1717) );
  NBUFFX2_RVT U2776 ( .A(n2918), .Y(n1699) );
  NBUFFX2_RVT U2777 ( .A(n2912), .Y(n1696) );
  NOR4X1_RVT U2778 ( .A1(n1854), .A2(n1853), .A3(n1852), .A4(n1851), .Y(n3006)
         );
  NBUFFX2_RVT U2779 ( .A(n1747), .Y(n1744) );
  NBUFFX2_RVT U2780 ( .A(n1737), .Y(n1735) );
  NBUFFX2_RVT U2781 ( .A(n1737), .Y(n1736) );
  NBUFFX2_RVT U2782 ( .A(n1723), .Y(n1718) );
  NBUFFX2_RVT U2783 ( .A(n1715), .Y(n1713) );
  NBUFFX2_RVT U2784 ( .A(n1715), .Y(n1714) );
  INVX1_RVT U2785 ( .A(search_data[30]), .Y(n1765) );
  INVX1_RVT U2786 ( .A(search_data[28]), .Y(n1759) );
  INVX1_RVT U2787 ( .A(n3007), .Y(n2989) );
  NOR4X1_RVT U2788 ( .A1(n1818), .A2(n1817), .A3(n1816), .A4(n1815), .Y(n3007)
         );
  NBUFFX2_RVT U2789 ( .A(n2942), .Y(n1742) );
  NBUFFX2_RVT U2790 ( .A(n1747), .Y(n1746) );
  NBUFFX2_RVT U2791 ( .A(n1737), .Y(n1734) );
  NBUFFX2_RVT U2792 ( .A(n2934), .Y(n1732) );
  NBUFFX2_RVT U2793 ( .A(n1729), .Y(n1727) );
  NBUFFX2_RVT U2794 ( .A(n2931), .Y(n1724) );
  NBUFFX2_RVT U2795 ( .A(n1723), .Y(n1719) );
  NBUFFX2_RVT U2796 ( .A(n2929), .Y(n1716) );
  NBUFFX2_RVT U2797 ( .A(n1723), .Y(n1722) );
  NBUFFX2_RVT U2798 ( .A(n1715), .Y(n1712) );
  NBUFFX2_RVT U2799 ( .A(n2923), .Y(n1710) );
  NBUFFX2_RVT U2800 ( .A(n1707), .Y(n1705) );
  NBUFFX2_RVT U2801 ( .A(n2920), .Y(n1701) );
  NBUFFX2_RVT U2802 ( .A(n2918), .Y(n1698) );
  NBUFFX2_RVT U2803 ( .A(n2912), .Y(n1695) );
  NBUFFX2_RVT U2804 ( .A(n1693), .Y(n1691) );
  INVX1_RVT U2805 ( .A(search_data[0]), .Y(n1751) );
  INVX1_RVT U2806 ( .A(search_data[0]), .Y(n1753) );
  AND2X1_RVT U2807 ( .A1(n3012), .A2(n2986), .Y(n1689) );
  NAND2X0_RVT U2808 ( .A1(n1771), .A2(n1769), .Y(n1782) );
  NAND2X0_RVT U2809 ( .A1(read_index[0]), .A2(n1769), .Y(n1780) );
  NAND2X0_RVT U2810 ( .A1(read_index[0]), .A2(read_index[1]), .Y(n1779) );
  AO22X1_RVT U2811 ( .A1(n1776), .A2(\words[9]/valid_o ), .A3(n1775), .A4(
        \words[11]/valid_o ), .Y(n1770) );
  NAND2X0_RVT U2812 ( .A1(read_index[1]), .A2(n1771), .Y(n1781) );
  AOI22X1_RVT U2813 ( .A1(n1776), .A2(\words[13]/valid_o ), .A3(n1775), .A4(
        \words[15]/valid_o ), .Y(n1773) );
  NAND2X0_RVT U2814 ( .A1(n1777), .A2(\words[12]/valid_o ), .Y(n1772) );
  AO22X1_RVT U2815 ( .A1(n1776), .A2(\words[1]/valid_o ), .A3(n1775), .A4(
        \words[3]/valid_o ), .Y(n1774) );
  AO22X1_RVT U2816 ( .A1(search_data[28]), .A2(\read_value_mux[0][28] ), .A3(
        n1757), .A4(n1636), .Y(n1783) );
  OA221X1_RVT U2817 ( .A1(search_data[1]), .A2(n11), .A3(n1754), .A4(
        \read_value_mux[0][1] ), .A5(n1783), .Y(n1790) );
  AO22X1_RVT U2818 ( .A1(search_data[30]), .A2(\read_value_mux[0][30] ), .A3(
        n1763), .A4(n12), .Y(n1784) );
  OA221X1_RVT U2819 ( .A1(search_data[29]), .A2(n1643), .A3(n1760), .A4(
        \read_value_mux[0][29] ), .A5(n1784), .Y(n1789) );
  AOI22X1_RVT U2820 ( .A1(n1543), .A2(\read_value_mux[0][26] ), .A3(n1542), 
        .A4(\read_value_mux[0][27] ), .Y(n1785) );
  OA221X1_RVT U2821 ( .A1(n1542), .A2(\read_value_mux[0][27] ), .A3(n1691), 
        .A4(\read_value_mux[0][26] ), .A5(n1785), .Y(n1788) );
  AOI22X1_RVT U2822 ( .A1(n1541), .A2(\read_value_mux[0][24] ), .A3(n1540), 
        .A4(\read_value_mux[0][25] ), .Y(n1786) );
  OA221X1_RVT U2823 ( .A1(n1540), .A2(\read_value_mux[0][25] ), .A3(n1695), 
        .A4(\read_value_mux[0][24] ), .A5(n1786), .Y(n1787) );
  NAND4X0_RVT U2824 ( .A1(n1790), .A2(n1789), .A3(n1788), .A4(n1787), .Y(n1818) );
  AOI22X1_RVT U2825 ( .A1(n1539), .A2(\read_value_mux[0][22] ), .A3(n1538), 
        .A4(\read_value_mux[0][23] ), .Y(n1791) );
  OA221X1_RVT U2826 ( .A1(n1538), .A2(\read_value_mux[0][23] ), .A3(n1698), 
        .A4(\read_value_mux[0][22] ), .A5(n1791), .Y(n1798) );
  AOI22X1_RVT U2827 ( .A1(n1537), .A2(\read_value_mux[0][20] ), .A3(n1536), 
        .A4(\read_value_mux[0][21] ), .Y(n1792) );
  OA221X1_RVT U2828 ( .A1(n1703), .A2(\read_value_mux[0][21] ), .A3(n1701), 
        .A4(\read_value_mux[0][20] ), .A5(n1792), .Y(n1797) );
  AOI22X1_RVT U2829 ( .A1(n1535), .A2(\read_value_mux[0][18] ), .A3(n1534), 
        .A4(\read_value_mux[0][19] ), .Y(n1793) );
  OA221X1_RVT U2830 ( .A1(n1708), .A2(\read_value_mux[0][19] ), .A3(n1705), 
        .A4(\read_value_mux[0][18] ), .A5(n1793), .Y(n1796) );
  AOI22X1_RVT U2831 ( .A1(n1533), .A2(\read_value_mux[0][16] ), .A3(n1712), 
        .A4(\read_value_mux[0][17] ), .Y(n1794) );
  OA221X1_RVT U2832 ( .A1(n1715), .A2(\read_value_mux[0][17] ), .A3(n1710), 
        .A4(\read_value_mux[0][16] ), .A5(n1794), .Y(n1795) );
  NAND4X0_RVT U2833 ( .A1(n1798), .A2(n1797), .A3(n1796), .A4(n1795), .Y(n1817) );
  AOI22X1_RVT U2834 ( .A1(n1532), .A2(\read_value_mux[0][14] ), .A3(n1719), 
        .A4(\read_value_mux[0][15] ), .Y(n1799) );
  OA221X1_RVT U2835 ( .A1(n1722), .A2(\read_value_mux[0][15] ), .A3(n1716), 
        .A4(\read_value_mux[0][14] ), .A5(n1799), .Y(n1806) );
  AOI22X1_RVT U2836 ( .A1(n1531), .A2(\read_value_mux[0][12] ), .A3(n1530), 
        .A4(\read_value_mux[0][13] ), .Y(n1800) );
  OA221X1_RVT U2837 ( .A1(n1530), .A2(\read_value_mux[0][13] ), .A3(n1724), 
        .A4(\read_value_mux[0][12] ), .A5(n1800), .Y(n1805) );
  AOI22X1_RVT U2838 ( .A1(n1529), .A2(\read_value_mux[0][10] ), .A3(n1528), 
        .A4(\read_value_mux[0][11] ), .Y(n1801) );
  OA221X1_RVT U2839 ( .A1(n1730), .A2(\read_value_mux[0][11] ), .A3(n1727), 
        .A4(\read_value_mux[0][10] ), .A5(n1801), .Y(n1804) );
  AOI22X1_RVT U2840 ( .A1(n1527), .A2(\read_value_mux[0][8] ), .A3(n1734), 
        .A4(\read_value_mux[0][9] ), .Y(n1802) );
  OA221X1_RVT U2841 ( .A1(n1737), .A2(\read_value_mux[0][9] ), .A3(n1732), 
        .A4(\read_value_mux[0][8] ), .A5(n1802), .Y(n1803) );
  NAND4X0_RVT U2842 ( .A1(n1806), .A2(n1805), .A3(n1804), .A4(n1803), .Y(n1816) );
  AOI22X1_RVT U2843 ( .A1(n2940), .A2(\read_value_mux[0][6] ), .A3(n1741), 
        .A4(\read_value_mux[0][7] ), .Y(n1807) );
  OA221X1_RVT U2844 ( .A1(n1739), .A2(\read_value_mux[0][7] ), .A3(n1738), 
        .A4(\read_value_mux[0][6] ), .A5(n1807), .Y(n1814) );
  AOI22X1_RVT U2845 ( .A1(n1526), .A2(\read_value_mux[0][4] ), .A3(n1525), 
        .A4(\read_value_mux[0][5] ), .Y(n1808) );
  OA221X1_RVT U2846 ( .A1(n1746), .A2(\read_value_mux[0][5] ), .A3(n1742), 
        .A4(\read_value_mux[0][4] ), .A5(n1808), .Y(n1813) );
  AOI22X1_RVT U2847 ( .A1(n1524), .A2(\read_value_mux[0][2] ), .A3(n1750), 
        .A4(\read_value_mux[0][3] ), .Y(n1809) );
  OA221X1_RVT U2848 ( .A1(n1750), .A2(\read_value_mux[0][3] ), .A3(n1524), 
        .A4(\read_value_mux[0][2] ), .A5(n1809), .Y(n1812) );
  OA221X1_RVT U2849 ( .A1(search_data[0]), .A2(n1644), .A3(n1751), .A4(
        \read_value_mux[0][0] ), .A5(search), .Y(n1810) );
  OA221X1_RVT U2850 ( .A1(search_data[31]), .A2(n1645), .A3(n1766), .A4(
        \read_value_mux[0][31] ), .A5(n1810), .Y(n1811) );
  NAND4X0_RVT U2851 ( .A1(n1814), .A2(n1813), .A3(n1812), .A4(n1811), .Y(n1815) );
  AO22X1_RVT U2852 ( .A1(search_data[28]), .A2(\read_value_mux[2][28] ), .A3(
        n1759), .A4(n1639), .Y(n1819) );
  OA221X1_RVT U2853 ( .A1(search_data[1]), .A2(n16), .A3(n1756), .A4(
        \read_value_mux[2][1] ), .A5(n1819), .Y(n1826) );
  AO22X1_RVT U2854 ( .A1(search_data[30]), .A2(\read_value_mux[2][30] ), .A3(
        n1765), .A4(n17), .Y(n1820) );
  OA221X1_RVT U2855 ( .A1(search_data[29]), .A2(n1658), .A3(n1762), .A4(
        \read_value_mux[2][29] ), .A5(n1820), .Y(n1825) );
  AOI22X1_RVT U2856 ( .A1(n1543), .A2(\read_value_mux[2][26] ), .A3(n1542), 
        .A4(\read_value_mux[2][27] ), .Y(n1821) );
  OA221X1_RVT U2857 ( .A1(n1542), .A2(\read_value_mux[2][27] ), .A3(n1691), 
        .A4(\read_value_mux[2][26] ), .A5(n1821), .Y(n1824) );
  AOI22X1_RVT U2858 ( .A1(n1541), .A2(\read_value_mux[2][24] ), .A3(n1540), 
        .A4(\read_value_mux[2][25] ), .Y(n1822) );
  OA221X1_RVT U2859 ( .A1(n1540), .A2(\read_value_mux[2][25] ), .A3(n1695), 
        .A4(\read_value_mux[2][24] ), .A5(n1822), .Y(n1823) );
  NAND4X0_RVT U2860 ( .A1(n1826), .A2(n1825), .A3(n1824), .A4(n1823), .Y(n1854) );
  AOI22X1_RVT U2861 ( .A1(n1539), .A2(\read_value_mux[2][22] ), .A3(n1538), 
        .A4(\read_value_mux[2][23] ), .Y(n1827) );
  OA221X1_RVT U2862 ( .A1(n1538), .A2(\read_value_mux[2][23] ), .A3(n1698), 
        .A4(\read_value_mux[2][22] ), .A5(n1827), .Y(n1834) );
  AOI22X1_RVT U2863 ( .A1(n1537), .A2(\read_value_mux[2][20] ), .A3(n1536), 
        .A4(\read_value_mux[2][21] ), .Y(n1828) );
  OA221X1_RVT U2864 ( .A1(n1703), .A2(\read_value_mux[2][21] ), .A3(n1701), 
        .A4(\read_value_mux[2][20] ), .A5(n1828), .Y(n1833) );
  AOI22X1_RVT U2865 ( .A1(n1535), .A2(\read_value_mux[2][18] ), .A3(n1534), 
        .A4(\read_value_mux[2][19] ), .Y(n1829) );
  OA221X1_RVT U2866 ( .A1(n1708), .A2(\read_value_mux[2][19] ), .A3(n1705), 
        .A4(\read_value_mux[2][18] ), .A5(n1829), .Y(n1832) );
  AOI22X1_RVT U2867 ( .A1(n1533), .A2(\read_value_mux[2][16] ), .A3(n1713), 
        .A4(\read_value_mux[2][17] ), .Y(n1830) );
  OA221X1_RVT U2868 ( .A1(n1714), .A2(\read_value_mux[2][17] ), .A3(n1710), 
        .A4(\read_value_mux[2][16] ), .A5(n1830), .Y(n1831) );
  NAND4X0_RVT U2869 ( .A1(n1834), .A2(n1833), .A3(n1832), .A4(n1831), .Y(n1853) );
  AOI22X1_RVT U2870 ( .A1(n1532), .A2(\read_value_mux[2][14] ), .A3(n1718), 
        .A4(\read_value_mux[2][15] ), .Y(n1835) );
  OA221X1_RVT U2871 ( .A1(n1722), .A2(\read_value_mux[2][15] ), .A3(n1716), 
        .A4(\read_value_mux[2][14] ), .A5(n1835), .Y(n1842) );
  AOI22X1_RVT U2872 ( .A1(n1531), .A2(\read_value_mux[2][12] ), .A3(n1530), 
        .A4(\read_value_mux[2][13] ), .Y(n1836) );
  OA221X1_RVT U2873 ( .A1(n1530), .A2(\read_value_mux[2][13] ), .A3(n1724), 
        .A4(\read_value_mux[2][12] ), .A5(n1836), .Y(n1841) );
  AOI22X1_RVT U2874 ( .A1(n1529), .A2(\read_value_mux[2][10] ), .A3(n1528), 
        .A4(\read_value_mux[2][11] ), .Y(n1837) );
  OA221X1_RVT U2875 ( .A1(n1730), .A2(\read_value_mux[2][11] ), .A3(n1727), 
        .A4(\read_value_mux[2][10] ), .A5(n1837), .Y(n1840) );
  AOI22X1_RVT U2876 ( .A1(n1527), .A2(\read_value_mux[2][8] ), .A3(n1735), 
        .A4(\read_value_mux[2][9] ), .Y(n1838) );
  OA221X1_RVT U2877 ( .A1(n1736), .A2(\read_value_mux[2][9] ), .A3(n1732), 
        .A4(\read_value_mux[2][8] ), .A5(n1838), .Y(n1839) );
  NAND4X0_RVT U2878 ( .A1(n1842), .A2(n1841), .A3(n1840), .A4(n1839), .Y(n1852) );
  AOI22X1_RVT U2879 ( .A1(n2940), .A2(\read_value_mux[2][6] ), .A3(n1741), 
        .A4(\read_value_mux[2][7] ), .Y(n1843) );
  OA221X1_RVT U2880 ( .A1(n1740), .A2(\read_value_mux[2][7] ), .A3(n1738), 
        .A4(\read_value_mux[2][6] ), .A5(n1843), .Y(n1850) );
  AOI22X1_RVT U2881 ( .A1(n1526), .A2(\read_value_mux[2][4] ), .A3(n1744), 
        .A4(\read_value_mux[2][5] ), .Y(n1844) );
  OA221X1_RVT U2882 ( .A1(n1746), .A2(\read_value_mux[2][5] ), .A3(n1742), 
        .A4(\read_value_mux[2][4] ), .A5(n1844), .Y(n1849) );
  AOI22X1_RVT U2883 ( .A1(n1524), .A2(\read_value_mux[2][2] ), .A3(n1750), 
        .A4(\read_value_mux[2][3] ), .Y(n1845) );
  OA221X1_RVT U2884 ( .A1(n1750), .A2(\read_value_mux[2][3] ), .A3(n1524), 
        .A4(\read_value_mux[2][2] ), .A5(n1845), .Y(n1848) );
  OA221X1_RVT U2885 ( .A1(search_data[0]), .A2(n1659), .A3(n1753), .A4(
        \read_value_mux[2][0] ), .A5(search), .Y(n1846) );
  OA221X1_RVT U2886 ( .A1(search_data[31]), .A2(n1660), .A3(n1768), .A4(
        \read_value_mux[2][31] ), .A5(n1846), .Y(n1847) );
  NAND4X0_RVT U2887 ( .A1(n1850), .A2(n1849), .A3(n1848), .A4(n1847), .Y(n1851) );
  AO22X1_RVT U2888 ( .A1(search_data[28]), .A2(\read_value_mux[3][28] ), .A3(
        n1759), .A4(n1637), .Y(n1855) );
  OA221X1_RVT U2889 ( .A1(search_data[1]), .A2(n18), .A3(n1756), .A4(
        \read_value_mux[3][1] ), .A5(n1855), .Y(n1862) );
  AO22X1_RVT U2890 ( .A1(search_data[30]), .A2(\read_value_mux[3][30] ), .A3(
        n1765), .A4(n19), .Y(n1856) );
  OA221X1_RVT U2891 ( .A1(search_data[29]), .A2(n1646), .A3(n1762), .A4(
        \read_value_mux[3][29] ), .A5(n1856), .Y(n1861) );
  AOI22X1_RVT U2892 ( .A1(n1691), .A2(\read_value_mux[3][26] ), .A3(n1542), 
        .A4(\read_value_mux[3][27] ), .Y(n1857) );
  OA221X1_RVT U2893 ( .A1(n1542), .A2(\read_value_mux[3][27] ), .A3(n1691), 
        .A4(\read_value_mux[3][26] ), .A5(n1857), .Y(n1860) );
  AOI22X1_RVT U2894 ( .A1(n1696), .A2(\read_value_mux[3][24] ), .A3(n1540), 
        .A4(\read_value_mux[3][25] ), .Y(n1858) );
  OA221X1_RVT U2895 ( .A1(n1540), .A2(\read_value_mux[3][25] ), .A3(n1695), 
        .A4(\read_value_mux[3][24] ), .A5(n1858), .Y(n1859) );
  NAND4X0_RVT U2896 ( .A1(n1862), .A2(n1861), .A3(n1860), .A4(n1859), .Y(n1890) );
  AOI22X1_RVT U2897 ( .A1(n1699), .A2(\read_value_mux[3][22] ), .A3(n1538), 
        .A4(\read_value_mux[3][23] ), .Y(n1863) );
  OA221X1_RVT U2898 ( .A1(n1538), .A2(\read_value_mux[3][23] ), .A3(n1698), 
        .A4(\read_value_mux[3][22] ), .A5(n1863), .Y(n1870) );
  AOI22X1_RVT U2899 ( .A1(n1537), .A2(\read_value_mux[3][20] ), .A3(n1536), 
        .A4(\read_value_mux[3][21] ), .Y(n1864) );
  OA221X1_RVT U2900 ( .A1(n1703), .A2(\read_value_mux[3][21] ), .A3(n1701), 
        .A4(\read_value_mux[3][20] ), .A5(n1864), .Y(n1869) );
  AOI22X1_RVT U2901 ( .A1(n1705), .A2(\read_value_mux[3][18] ), .A3(n1534), 
        .A4(\read_value_mux[3][19] ), .Y(n1865) );
  OA221X1_RVT U2902 ( .A1(n1708), .A2(\read_value_mux[3][19] ), .A3(n1705), 
        .A4(\read_value_mux[3][18] ), .A5(n1865), .Y(n1868) );
  AOI22X1_RVT U2903 ( .A1(n1533), .A2(\read_value_mux[3][16] ), .A3(n1712), 
        .A4(\read_value_mux[3][17] ), .Y(n1866) );
  OA221X1_RVT U2904 ( .A1(n1714), .A2(\read_value_mux[3][17] ), .A3(n1710), 
        .A4(\read_value_mux[3][16] ), .A5(n1866), .Y(n1867) );
  NAND4X0_RVT U2905 ( .A1(n1870), .A2(n1869), .A3(n1868), .A4(n1867), .Y(n1889) );
  AOI22X1_RVT U2906 ( .A1(n1717), .A2(\read_value_mux[3][14] ), .A3(n1718), 
        .A4(\read_value_mux[3][15] ), .Y(n1871) );
  OA221X1_RVT U2907 ( .A1(n1722), .A2(\read_value_mux[3][15] ), .A3(n1716), 
        .A4(\read_value_mux[3][14] ), .A5(n1871), .Y(n1878) );
  AOI22X1_RVT U2908 ( .A1(n1725), .A2(\read_value_mux[3][12] ), .A3(n1530), 
        .A4(\read_value_mux[3][13] ), .Y(n1872) );
  OA221X1_RVT U2909 ( .A1(n1530), .A2(\read_value_mux[3][13] ), .A3(n1724), 
        .A4(\read_value_mux[3][12] ), .A5(n1872), .Y(n1877) );
  AOI22X1_RVT U2910 ( .A1(n1727), .A2(\read_value_mux[3][10] ), .A3(n1528), 
        .A4(\read_value_mux[3][11] ), .Y(n1873) );
  OA221X1_RVT U2911 ( .A1(n1730), .A2(\read_value_mux[3][11] ), .A3(n1727), 
        .A4(\read_value_mux[3][10] ), .A5(n1873), .Y(n1876) );
  AOI22X1_RVT U2912 ( .A1(n1733), .A2(\read_value_mux[3][8] ), .A3(n1734), 
        .A4(\read_value_mux[3][9] ), .Y(n1874) );
  OA221X1_RVT U2913 ( .A1(n1736), .A2(\read_value_mux[3][9] ), .A3(n1732), 
        .A4(\read_value_mux[3][8] ), .A5(n1874), .Y(n1875) );
  NAND4X0_RVT U2914 ( .A1(n1878), .A2(n1877), .A3(n1876), .A4(n1875), .Y(n1888) );
  AOI22X1_RVT U2915 ( .A1(n1738), .A2(\read_value_mux[3][6] ), .A3(n1741), 
        .A4(\read_value_mux[3][7] ), .Y(n1879) );
  OA221X1_RVT U2916 ( .A1(n1739), .A2(\read_value_mux[3][7] ), .A3(n1738), 
        .A4(\read_value_mux[3][6] ), .A5(n1879), .Y(n1886) );
  AOI22X1_RVT U2917 ( .A1(n1743), .A2(\read_value_mux[3][4] ), .A3(n1744), 
        .A4(\read_value_mux[3][5] ), .Y(n1880) );
  OA221X1_RVT U2918 ( .A1(n1746), .A2(\read_value_mux[3][5] ), .A3(n1742), 
        .A4(\read_value_mux[3][4] ), .A5(n1880), .Y(n1885) );
  AOI22X1_RVT U2919 ( .A1(n1748), .A2(\read_value_mux[3][2] ), .A3(n1750), 
        .A4(\read_value_mux[3][3] ), .Y(n1881) );
  OA221X1_RVT U2920 ( .A1(n1750), .A2(\read_value_mux[3][3] ), .A3(n1524), 
        .A4(\read_value_mux[3][2] ), .A5(n1881), .Y(n1884) );
  OA221X1_RVT U2921 ( .A1(search_data[0]), .A2(n1647), .A3(n1753), .A4(
        \read_value_mux[3][0] ), .A5(search), .Y(n1882) );
  OA221X1_RVT U2922 ( .A1(search_data[31]), .A2(n1648), .A3(n1768), .A4(
        \read_value_mux[3][31] ), .A5(n1882), .Y(n1883) );
  NAND4X0_RVT U2923 ( .A1(n1886), .A2(n1885), .A3(n1884), .A4(n1883), .Y(n1887) );
  AO22X1_RVT U2924 ( .A1(search_data[28]), .A2(\read_value_mux[5][28] ), .A3(
        n1759), .A4(n1557), .Y(n1891) );
  OA221X1_RVT U2925 ( .A1(search_data[1]), .A2(n23), .A3(n1756), .A4(
        \read_value_mux[5][1] ), .A5(n1891), .Y(n1898) );
  AO22X1_RVT U2926 ( .A1(search_data[30]), .A2(\read_value_mux[5][30] ), .A3(
        n1765), .A4(n24), .Y(n1892) );
  OA221X1_RVT U2927 ( .A1(search_data[29]), .A2(n1661), .A3(n1762), .A4(
        \read_value_mux[5][29] ), .A5(n1892), .Y(n1897) );
  AOI22X1_RVT U2928 ( .A1(n1692), .A2(\read_value_mux[5][26] ), .A3(n1542), 
        .A4(\read_value_mux[5][27] ), .Y(n1893) );
  OA221X1_RVT U2929 ( .A1(n1542), .A2(\read_value_mux[5][27] ), .A3(n1692), 
        .A4(\read_value_mux[5][26] ), .A5(n1893), .Y(n1896) );
  AOI22X1_RVT U2930 ( .A1(n1696), .A2(\read_value_mux[5][24] ), .A3(n1540), 
        .A4(\read_value_mux[5][25] ), .Y(n1894) );
  OA221X1_RVT U2931 ( .A1(n1540), .A2(\read_value_mux[5][25] ), .A3(n1696), 
        .A4(\read_value_mux[5][24] ), .A5(n1894), .Y(n1895) );
  NAND4X0_RVT U2932 ( .A1(n1898), .A2(n1897), .A3(n1896), .A4(n1895), .Y(n1926) );
  AOI22X1_RVT U2933 ( .A1(n1699), .A2(\read_value_mux[5][22] ), .A3(n1538), 
        .A4(\read_value_mux[5][23] ), .Y(n1899) );
  OA221X1_RVT U2934 ( .A1(n1538), .A2(\read_value_mux[5][23] ), .A3(n1699), 
        .A4(\read_value_mux[5][22] ), .A5(n1899), .Y(n1906) );
  AOI22X1_RVT U2935 ( .A1(n1702), .A2(\read_value_mux[5][20] ), .A3(n1703), 
        .A4(\read_value_mux[5][21] ), .Y(n1900) );
  OA221X1_RVT U2936 ( .A1(n1703), .A2(\read_value_mux[5][21] ), .A3(n1702), 
        .A4(\read_value_mux[5][20] ), .A5(n1900), .Y(n1905) );
  AOI22X1_RVT U2937 ( .A1(n1706), .A2(\read_value_mux[5][18] ), .A3(n1708), 
        .A4(\read_value_mux[5][19] ), .Y(n1901) );
  OA221X1_RVT U2938 ( .A1(n1708), .A2(\read_value_mux[5][19] ), .A3(n1706), 
        .A4(\read_value_mux[5][18] ), .A5(n1901), .Y(n1904) );
  AOI22X1_RVT U2939 ( .A1(n1711), .A2(\read_value_mux[5][16] ), .A3(n1713), 
        .A4(\read_value_mux[5][17] ), .Y(n1902) );
  OA221X1_RVT U2940 ( .A1(n1714), .A2(\read_value_mux[5][17] ), .A3(n1711), 
        .A4(\read_value_mux[5][16] ), .A5(n1902), .Y(n1903) );
  NAND4X0_RVT U2941 ( .A1(n1906), .A2(n1905), .A3(n1904), .A4(n1903), .Y(n1925) );
  AOI22X1_RVT U2942 ( .A1(n1717), .A2(\read_value_mux[5][14] ), .A3(n1718), 
        .A4(\read_value_mux[5][15] ), .Y(n1907) );
  OA221X1_RVT U2943 ( .A1(n1722), .A2(\read_value_mux[5][15] ), .A3(n1717), 
        .A4(\read_value_mux[5][14] ), .A5(n1907), .Y(n1914) );
  AOI22X1_RVT U2944 ( .A1(n1725), .A2(\read_value_mux[5][12] ), .A3(n1530), 
        .A4(\read_value_mux[5][13] ), .Y(n1908) );
  OA221X1_RVT U2945 ( .A1(n1530), .A2(\read_value_mux[5][13] ), .A3(n1725), 
        .A4(\read_value_mux[5][12] ), .A5(n1908), .Y(n1913) );
  AOI22X1_RVT U2946 ( .A1(n1728), .A2(\read_value_mux[5][10] ), .A3(n1730), 
        .A4(\read_value_mux[5][11] ), .Y(n1909) );
  OA221X1_RVT U2947 ( .A1(n1730), .A2(\read_value_mux[5][11] ), .A3(n1728), 
        .A4(\read_value_mux[5][10] ), .A5(n1909), .Y(n1912) );
  AOI22X1_RVT U2948 ( .A1(n1733), .A2(\read_value_mux[5][8] ), .A3(n1735), 
        .A4(\read_value_mux[5][9] ), .Y(n1910) );
  OA221X1_RVT U2949 ( .A1(n1736), .A2(\read_value_mux[5][9] ), .A3(n1733), 
        .A4(\read_value_mux[5][8] ), .A5(n1910), .Y(n1911) );
  NAND4X0_RVT U2950 ( .A1(n1914), .A2(n1913), .A3(n1912), .A4(n1911), .Y(n1924) );
  AOI22X1_RVT U2951 ( .A1(n1738), .A2(\read_value_mux[5][6] ), .A3(n1741), 
        .A4(\read_value_mux[5][7] ), .Y(n1915) );
  OA221X1_RVT U2952 ( .A1(n1739), .A2(\read_value_mux[5][7] ), .A3(n1738), 
        .A4(\read_value_mux[5][6] ), .A5(n1915), .Y(n1922) );
  AOI22X1_RVT U2953 ( .A1(n1743), .A2(\read_value_mux[5][4] ), .A3(n1744), 
        .A4(\read_value_mux[5][5] ), .Y(n1916) );
  OA221X1_RVT U2954 ( .A1(n1746), .A2(\read_value_mux[5][5] ), .A3(n1743), 
        .A4(\read_value_mux[5][4] ), .A5(n1916), .Y(n1921) );
  AOI22X1_RVT U2955 ( .A1(n1748), .A2(\read_value_mux[5][2] ), .A3(n1750), 
        .A4(\read_value_mux[5][3] ), .Y(n1917) );
  OA221X1_RVT U2956 ( .A1(n1750), .A2(\read_value_mux[5][3] ), .A3(n1748), 
        .A4(\read_value_mux[5][2] ), .A5(n1917), .Y(n1920) );
  OA221X1_RVT U2957 ( .A1(search_data[0]), .A2(n1601), .A3(n1753), .A4(
        \read_value_mux[5][0] ), .A5(search), .Y(n1918) );
  OA221X1_RVT U2958 ( .A1(search_data[31]), .A2(n1662), .A3(n1768), .A4(
        \read_value_mux[5][31] ), .A5(n1918), .Y(n1919) );
  NAND4X0_RVT U2959 ( .A1(n1922), .A2(n1921), .A3(n1920), .A4(n1919), .Y(n1923) );
  AO22X1_RVT U2960 ( .A1(search_data[28]), .A2(\read_value_mux[7][28] ), .A3(
        n1759), .A4(n1544), .Y(n1927) );
  OA221X1_RVT U2961 ( .A1(search_data[1]), .A2(n28), .A3(n1756), .A4(
        \read_value_mux[7][1] ), .A5(n1927), .Y(n1934) );
  AO22X1_RVT U2962 ( .A1(search_data[30]), .A2(\read_value_mux[7][30] ), .A3(
        n1765), .A4(n29), .Y(n1928) );
  OA221X1_RVT U2963 ( .A1(search_data[29]), .A2(n1649), .A3(n1762), .A4(
        \read_value_mux[7][29] ), .A5(n1928), .Y(n1933) );
  AOI22X1_RVT U2964 ( .A1(n1543), .A2(\read_value_mux[7][26] ), .A3(n1694), 
        .A4(\read_value_mux[7][27] ), .Y(n1929) );
  OA221X1_RVT U2965 ( .A1(n1542), .A2(\read_value_mux[7][27] ), .A3(n1692), 
        .A4(\read_value_mux[7][26] ), .A5(n1929), .Y(n1932) );
  AOI22X1_RVT U2966 ( .A1(n1541), .A2(\read_value_mux[7][24] ), .A3(n1540), 
        .A4(\read_value_mux[7][25] ), .Y(n1930) );
  OA221X1_RVT U2967 ( .A1(n1540), .A2(\read_value_mux[7][25] ), .A3(n1696), 
        .A4(\read_value_mux[7][24] ), .A5(n1930), .Y(n1931) );
  NAND4X0_RVT U2968 ( .A1(n1934), .A2(n1933), .A3(n1932), .A4(n1931), .Y(n1962) );
  AOI22X1_RVT U2969 ( .A1(n1539), .A2(\read_value_mux[7][22] ), .A3(n1700), 
        .A4(\read_value_mux[7][23] ), .Y(n1935) );
  OA221X1_RVT U2970 ( .A1(n1538), .A2(\read_value_mux[7][23] ), .A3(n1699), 
        .A4(\read_value_mux[7][22] ), .A5(n1935), .Y(n1942) );
  AOI22X1_RVT U2971 ( .A1(n1537), .A2(\read_value_mux[7][20] ), .A3(n1536), 
        .A4(\read_value_mux[7][21] ), .Y(n1936) );
  OA221X1_RVT U2972 ( .A1(n1703), .A2(\read_value_mux[7][21] ), .A3(n1702), 
        .A4(\read_value_mux[7][20] ), .A5(n1936), .Y(n1941) );
  AOI22X1_RVT U2973 ( .A1(n1535), .A2(\read_value_mux[7][18] ), .A3(n1534), 
        .A4(\read_value_mux[7][19] ), .Y(n1937) );
  OA221X1_RVT U2974 ( .A1(n1708), .A2(\read_value_mux[7][19] ), .A3(n1706), 
        .A4(\read_value_mux[7][18] ), .A5(n1937), .Y(n1940) );
  AOI22X1_RVT U2975 ( .A1(n1533), .A2(\read_value_mux[7][16] ), .A3(n1712), 
        .A4(\read_value_mux[7][17] ), .Y(n1938) );
  OA221X1_RVT U2976 ( .A1(n1714), .A2(\read_value_mux[7][17] ), .A3(n1711), 
        .A4(\read_value_mux[7][16] ), .A5(n1938), .Y(n1939) );
  NAND4X0_RVT U2977 ( .A1(n1942), .A2(n1941), .A3(n1940), .A4(n1939), .Y(n1961) );
  AOI22X1_RVT U2978 ( .A1(n1532), .A2(\read_value_mux[7][14] ), .A3(n1718), 
        .A4(\read_value_mux[7][15] ), .Y(n1943) );
  OA221X1_RVT U2979 ( .A1(n1722), .A2(\read_value_mux[7][15] ), .A3(n1717), 
        .A4(\read_value_mux[7][14] ), .A5(n1943), .Y(n1950) );
  AOI22X1_RVT U2980 ( .A1(n1531), .A2(\read_value_mux[7][12] ), .A3(n1726), 
        .A4(\read_value_mux[7][13] ), .Y(n1944) );
  OA221X1_RVT U2981 ( .A1(n1530), .A2(\read_value_mux[7][13] ), .A3(n1725), 
        .A4(\read_value_mux[7][12] ), .A5(n1944), .Y(n1949) );
  AOI22X1_RVT U2982 ( .A1(n1529), .A2(\read_value_mux[7][10] ), .A3(n1528), 
        .A4(\read_value_mux[7][11] ), .Y(n1945) );
  OA221X1_RVT U2983 ( .A1(n1730), .A2(\read_value_mux[7][11] ), .A3(n1728), 
        .A4(\read_value_mux[7][10] ), .A5(n1945), .Y(n1948) );
  AOI22X1_RVT U2984 ( .A1(n1527), .A2(\read_value_mux[7][8] ), .A3(n1734), 
        .A4(\read_value_mux[7][9] ), .Y(n1946) );
  OA221X1_RVT U2985 ( .A1(n1736), .A2(\read_value_mux[7][9] ), .A3(n1733), 
        .A4(\read_value_mux[7][8] ), .A5(n1946), .Y(n1947) );
  NAND4X0_RVT U2986 ( .A1(n1950), .A2(n1949), .A3(n1948), .A4(n1947), .Y(n1960) );
  AOI22X1_RVT U2987 ( .A1(n2940), .A2(\read_value_mux[7][6] ), .A3(n1741), 
        .A4(\read_value_mux[7][7] ), .Y(n1951) );
  OA221X1_RVT U2988 ( .A1(n1739), .A2(\read_value_mux[7][7] ), .A3(n1738), 
        .A4(\read_value_mux[7][6] ), .A5(n1951), .Y(n1958) );
  AOI22X1_RVT U2989 ( .A1(n1526), .A2(\read_value_mux[7][4] ), .A3(n1744), 
        .A4(\read_value_mux[7][5] ), .Y(n1952) );
  OA221X1_RVT U2990 ( .A1(n1746), .A2(\read_value_mux[7][5] ), .A3(n1743), 
        .A4(\read_value_mux[7][4] ), .A5(n1952), .Y(n1957) );
  AOI22X1_RVT U2991 ( .A1(n1524), .A2(\read_value_mux[7][2] ), .A3(n1750), 
        .A4(\read_value_mux[7][3] ), .Y(n1953) );
  OA221X1_RVT U2992 ( .A1(n1750), .A2(\read_value_mux[7][3] ), .A3(n1748), 
        .A4(\read_value_mux[7][2] ), .A5(n1953), .Y(n1956) );
  OA221X1_RVT U2993 ( .A1(search_data[0]), .A2(n1568), .A3(n1753), .A4(
        \read_value_mux[7][0] ), .A5(search), .Y(n1954) );
  OA221X1_RVT U2994 ( .A1(search_data[31]), .A2(n1650), .A3(n1768), .A4(
        \read_value_mux[7][31] ), .A5(n1954), .Y(n1955) );
  NAND4X0_RVT U2995 ( .A1(n1958), .A2(n1957), .A3(n1956), .A4(n1955), .Y(n1959) );
  AO22X1_RVT U2996 ( .A1(search_data[28]), .A2(\read_value_mux[6][28] ), .A3(
        n1759), .A4(n1640), .Y(n1963) );
  OA221X1_RVT U2997 ( .A1(search_data[1]), .A2(n26), .A3(n1756), .A4(
        \read_value_mux[6][1] ), .A5(n1963), .Y(n1970) );
  AO22X1_RVT U2998 ( .A1(search_data[30]), .A2(\read_value_mux[6][30] ), .A3(
        n1765), .A4(n27), .Y(n1964) );
  OA221X1_RVT U2999 ( .A1(search_data[29]), .A2(n1663), .A3(n1762), .A4(
        \read_value_mux[6][29] ), .A5(n1964), .Y(n1969) );
  AOI22X1_RVT U3000 ( .A1(n1692), .A2(\read_value_mux[6][26] ), .A3(n1542), 
        .A4(\read_value_mux[6][27] ), .Y(n1965) );
  OA221X1_RVT U3001 ( .A1(n1542), .A2(\read_value_mux[6][27] ), .A3(n1692), 
        .A4(\read_value_mux[6][26] ), .A5(n1965), .Y(n1968) );
  AOI22X1_RVT U3002 ( .A1(n1696), .A2(\read_value_mux[6][24] ), .A3(n1697), 
        .A4(\read_value_mux[6][25] ), .Y(n1966) );
  OA221X1_RVT U3003 ( .A1(n1540), .A2(\read_value_mux[6][25] ), .A3(n1696), 
        .A4(\read_value_mux[6][24] ), .A5(n1966), .Y(n1967) );
  NAND4X0_RVT U3004 ( .A1(n1970), .A2(n1969), .A3(n1968), .A4(n1967), .Y(n1998) );
  AOI22X1_RVT U3005 ( .A1(n1699), .A2(\read_value_mux[6][22] ), .A3(n1538), 
        .A4(\read_value_mux[6][23] ), .Y(n1971) );
  OA221X1_RVT U3006 ( .A1(n1538), .A2(\read_value_mux[6][23] ), .A3(n1699), 
        .A4(\read_value_mux[6][22] ), .A5(n1971), .Y(n1978) );
  AOI22X1_RVT U3007 ( .A1(n1702), .A2(\read_value_mux[6][20] ), .A3(n1536), 
        .A4(\read_value_mux[6][21] ), .Y(n1972) );
  OA221X1_RVT U3008 ( .A1(n1703), .A2(\read_value_mux[6][21] ), .A3(n1702), 
        .A4(\read_value_mux[6][20] ), .A5(n1972), .Y(n1977) );
  AOI22X1_RVT U3009 ( .A1(n1706), .A2(\read_value_mux[6][18] ), .A3(n1534), 
        .A4(\read_value_mux[6][19] ), .Y(n1973) );
  OA221X1_RVT U3010 ( .A1(n1708), .A2(\read_value_mux[6][19] ), .A3(n1706), 
        .A4(\read_value_mux[6][18] ), .A5(n1973), .Y(n1976) );
  AOI22X1_RVT U3011 ( .A1(n1711), .A2(\read_value_mux[6][16] ), .A3(n1712), 
        .A4(\read_value_mux[6][17] ), .Y(n1974) );
  OA221X1_RVT U3012 ( .A1(n1714), .A2(\read_value_mux[6][17] ), .A3(n1711), 
        .A4(\read_value_mux[6][16] ), .A5(n1974), .Y(n1975) );
  NAND4X0_RVT U3013 ( .A1(n1978), .A2(n1977), .A3(n1976), .A4(n1975), .Y(n1997) );
  AOI22X1_RVT U3014 ( .A1(n1717), .A2(\read_value_mux[6][14] ), .A3(n1718), 
        .A4(\read_value_mux[6][15] ), .Y(n1979) );
  OA221X1_RVT U3015 ( .A1(n1722), .A2(\read_value_mux[6][15] ), .A3(n1717), 
        .A4(\read_value_mux[6][14] ), .A5(n1979), .Y(n1986) );
  AOI22X1_RVT U3016 ( .A1(n1725), .A2(\read_value_mux[6][12] ), .A3(n1530), 
        .A4(\read_value_mux[6][13] ), .Y(n1980) );
  OA221X1_RVT U3017 ( .A1(n1530), .A2(\read_value_mux[6][13] ), .A3(n1725), 
        .A4(\read_value_mux[6][12] ), .A5(n1980), .Y(n1985) );
  AOI22X1_RVT U3018 ( .A1(n1728), .A2(\read_value_mux[6][10] ), .A3(n1528), 
        .A4(\read_value_mux[6][11] ), .Y(n1981) );
  OA221X1_RVT U3019 ( .A1(n1730), .A2(\read_value_mux[6][11] ), .A3(n1728), 
        .A4(\read_value_mux[6][10] ), .A5(n1981), .Y(n1984) );
  AOI22X1_RVT U3020 ( .A1(n1733), .A2(\read_value_mux[6][8] ), .A3(n1734), 
        .A4(\read_value_mux[6][9] ), .Y(n1982) );
  OA221X1_RVT U3021 ( .A1(n1736), .A2(\read_value_mux[6][9] ), .A3(n1733), 
        .A4(\read_value_mux[6][8] ), .A5(n1982), .Y(n1983) );
  NAND4X0_RVT U3022 ( .A1(n1986), .A2(n1985), .A3(n1984), .A4(n1983), .Y(n1996) );
  AOI22X1_RVT U3023 ( .A1(n1738), .A2(\read_value_mux[6][6] ), .A3(n1741), 
        .A4(\read_value_mux[6][7] ), .Y(n1987) );
  OA221X1_RVT U3024 ( .A1(n1739), .A2(\read_value_mux[6][7] ), .A3(n1738), 
        .A4(\read_value_mux[6][6] ), .A5(n1987), .Y(n1994) );
  AOI22X1_RVT U3025 ( .A1(n1743), .A2(\read_value_mux[6][4] ), .A3(n1744), 
        .A4(\read_value_mux[6][5] ), .Y(n1988) );
  OA221X1_RVT U3026 ( .A1(n1746), .A2(\read_value_mux[6][5] ), .A3(n1743), 
        .A4(\read_value_mux[6][4] ), .A5(n1988), .Y(n1993) );
  AOI22X1_RVT U3027 ( .A1(n1748), .A2(\read_value_mux[6][2] ), .A3(n1750), 
        .A4(\read_value_mux[6][3] ), .Y(n1989) );
  OA221X1_RVT U3028 ( .A1(n1750), .A2(\read_value_mux[6][3] ), .A3(n1748), 
        .A4(\read_value_mux[6][2] ), .A5(n1989), .Y(n1992) );
  OA221X1_RVT U3029 ( .A1(search_data[0]), .A2(n1664), .A3(n1753), .A4(
        \read_value_mux[6][0] ), .A5(search), .Y(n1990) );
  OA221X1_RVT U3030 ( .A1(search_data[31]), .A2(n1665), .A3(n1768), .A4(
        \read_value_mux[6][31] ), .A5(n1990), .Y(n1991) );
  NAND4X0_RVT U3031 ( .A1(n1994), .A2(n1993), .A3(n1992), .A4(n1991), .Y(n1995) );
  AO22X1_RVT U3032 ( .A1(search_data[28]), .A2(\read_value_mux[4][28] ), .A3(
        n1759), .A4(n1638), .Y(n1999) );
  OA221X1_RVT U3033 ( .A1(search_data[1]), .A2(n21), .A3(n1756), .A4(
        \read_value_mux[4][1] ), .A5(n1999), .Y(n2006) );
  AO22X1_RVT U3034 ( .A1(search_data[30]), .A2(\read_value_mux[4][30] ), .A3(
        n1765), .A4(n22), .Y(n2000) );
  OA221X1_RVT U3035 ( .A1(search_data[29]), .A2(n1651), .A3(n1762), .A4(
        \read_value_mux[4][29] ), .A5(n2000), .Y(n2005) );
  AOI22X1_RVT U3036 ( .A1(n1543), .A2(\read_value_mux[4][26] ), .A3(n1542), 
        .A4(\read_value_mux[4][27] ), .Y(n2001) );
  OA221X1_RVT U3037 ( .A1(n1542), .A2(\read_value_mux[4][27] ), .A3(n1691), 
        .A4(\read_value_mux[4][26] ), .A5(n2001), .Y(n2004) );
  AOI22X1_RVT U3038 ( .A1(n1541), .A2(\read_value_mux[4][24] ), .A3(n1540), 
        .A4(\read_value_mux[4][25] ), .Y(n2002) );
  OA221X1_RVT U3039 ( .A1(n1540), .A2(\read_value_mux[4][25] ), .A3(n1695), 
        .A4(\read_value_mux[4][24] ), .A5(n2002), .Y(n2003) );
  NAND4X0_RVT U3040 ( .A1(n2006), .A2(n2005), .A3(n2004), .A4(n2003), .Y(n2034) );
  AOI22X1_RVT U3041 ( .A1(n1539), .A2(\read_value_mux[4][22] ), .A3(n1538), 
        .A4(\read_value_mux[4][23] ), .Y(n2007) );
  OA221X1_RVT U3042 ( .A1(n1538), .A2(\read_value_mux[4][23] ), .A3(n1698), 
        .A4(\read_value_mux[4][22] ), .A5(n2007), .Y(n2014) );
  AOI22X1_RVT U3043 ( .A1(n1537), .A2(\read_value_mux[4][20] ), .A3(n1536), 
        .A4(\read_value_mux[4][21] ), .Y(n2008) );
  OA221X1_RVT U3044 ( .A1(n1703), .A2(\read_value_mux[4][21] ), .A3(n1701), 
        .A4(\read_value_mux[4][20] ), .A5(n2008), .Y(n2013) );
  AOI22X1_RVT U3045 ( .A1(n1535), .A2(\read_value_mux[4][18] ), .A3(n1534), 
        .A4(\read_value_mux[4][19] ), .Y(n2009) );
  OA221X1_RVT U3046 ( .A1(n1708), .A2(\read_value_mux[4][19] ), .A3(n1705), 
        .A4(\read_value_mux[4][18] ), .A5(n2009), .Y(n2012) );
  AOI22X1_RVT U3047 ( .A1(n1533), .A2(\read_value_mux[4][16] ), .A3(n1714), 
        .A4(\read_value_mux[4][17] ), .Y(n2010) );
  OA221X1_RVT U3048 ( .A1(n1714), .A2(\read_value_mux[4][17] ), .A3(n1710), 
        .A4(\read_value_mux[4][16] ), .A5(n2010), .Y(n2011) );
  NAND4X0_RVT U3049 ( .A1(n2014), .A2(n2013), .A3(n2012), .A4(n2011), .Y(n2033) );
  AOI22X1_RVT U3050 ( .A1(n1532), .A2(\read_value_mux[4][14] ), .A3(n1718), 
        .A4(\read_value_mux[4][15] ), .Y(n2015) );
  OA221X1_RVT U3051 ( .A1(n1722), .A2(\read_value_mux[4][15] ), .A3(n1716), 
        .A4(\read_value_mux[4][14] ), .A5(n2015), .Y(n2022) );
  AOI22X1_RVT U3052 ( .A1(n1531), .A2(\read_value_mux[4][12] ), .A3(n1530), 
        .A4(\read_value_mux[4][13] ), .Y(n2016) );
  OA221X1_RVT U3053 ( .A1(n1530), .A2(\read_value_mux[4][13] ), .A3(n1724), 
        .A4(\read_value_mux[4][12] ), .A5(n2016), .Y(n2021) );
  AOI22X1_RVT U3054 ( .A1(n1529), .A2(\read_value_mux[4][10] ), .A3(n1528), 
        .A4(\read_value_mux[4][11] ), .Y(n2017) );
  OA221X1_RVT U3055 ( .A1(n1730), .A2(\read_value_mux[4][11] ), .A3(n1727), 
        .A4(\read_value_mux[4][10] ), .A5(n2017), .Y(n2020) );
  AOI22X1_RVT U3056 ( .A1(n1527), .A2(\read_value_mux[4][8] ), .A3(n1736), 
        .A4(\read_value_mux[4][9] ), .Y(n2018) );
  OA221X1_RVT U3057 ( .A1(n1736), .A2(\read_value_mux[4][9] ), .A3(n1732), 
        .A4(\read_value_mux[4][8] ), .A5(n2018), .Y(n2019) );
  NAND4X0_RVT U3058 ( .A1(n2022), .A2(n2021), .A3(n2020), .A4(n2019), .Y(n2032) );
  AOI22X1_RVT U3059 ( .A1(n2940), .A2(\read_value_mux[4][6] ), .A3(n1741), 
        .A4(\read_value_mux[4][7] ), .Y(n2023) );
  OA221X1_RVT U3060 ( .A1(n1740), .A2(\read_value_mux[4][7] ), .A3(n1738), 
        .A4(\read_value_mux[4][6] ), .A5(n2023), .Y(n2030) );
  AOI22X1_RVT U3061 ( .A1(n1526), .A2(\read_value_mux[4][4] ), .A3(n1744), 
        .A4(\read_value_mux[4][5] ), .Y(n2024) );
  OA221X1_RVT U3062 ( .A1(n1746), .A2(\read_value_mux[4][5] ), .A3(n1742), 
        .A4(\read_value_mux[4][4] ), .A5(n2024), .Y(n2029) );
  AOI22X1_RVT U3063 ( .A1(n1524), .A2(\read_value_mux[4][2] ), .A3(n1750), 
        .A4(\read_value_mux[4][3] ), .Y(n2025) );
  OA221X1_RVT U3064 ( .A1(n1750), .A2(\read_value_mux[4][3] ), .A3(n1524), 
        .A4(\read_value_mux[4][2] ), .A5(n2025), .Y(n2028) );
  OA221X1_RVT U3065 ( .A1(search_data[0]), .A2(n1652), .A3(n1753), .A4(
        \read_value_mux[4][0] ), .A5(search), .Y(n2026) );
  OA221X1_RVT U3066 ( .A1(search_data[31]), .A2(n1653), .A3(n1768), .A4(
        \read_value_mux[4][31] ), .A5(n2026), .Y(n2027) );
  NAND4X0_RVT U3067 ( .A1(n2030), .A2(n2029), .A3(n2028), .A4(n2027), .Y(n2031) );
  AO22X1_RVT U3068 ( .A1(search_data[28]), .A2(\read_value_mux[1][28] ), .A3(
        n1758), .A4(n1641), .Y(n2035) );
  OA221X1_RVT U3069 ( .A1(search_data[1]), .A2(n14), .A3(n1755), .A4(
        \read_value_mux[1][1] ), .A5(n2035), .Y(n2042) );
  AO22X1_RVT U3070 ( .A1(search_data[30]), .A2(\read_value_mux[1][30] ), .A3(
        n1764), .A4(n15), .Y(n2036) );
  OA221X1_RVT U3071 ( .A1(search_data[29]), .A2(n1666), .A3(n1762), .A4(
        \read_value_mux[1][29] ), .A5(n2036), .Y(n2041) );
  AOI22X1_RVT U3072 ( .A1(n1692), .A2(\read_value_mux[1][26] ), .A3(n1542), 
        .A4(\read_value_mux[1][27] ), .Y(n2037) );
  OA221X1_RVT U3073 ( .A1(n1542), .A2(\read_value_mux[1][27] ), .A3(n1692), 
        .A4(\read_value_mux[1][26] ), .A5(n2037), .Y(n2040) );
  AOI22X1_RVT U3074 ( .A1(n1695), .A2(\read_value_mux[1][24] ), .A3(n1540), 
        .A4(\read_value_mux[1][25] ), .Y(n2038) );
  OA221X1_RVT U3075 ( .A1(n1540), .A2(\read_value_mux[1][25] ), .A3(n1696), 
        .A4(\read_value_mux[1][24] ), .A5(n2038), .Y(n2039) );
  NAND4X0_RVT U3076 ( .A1(n2042), .A2(n2041), .A3(n2040), .A4(n2039), .Y(n2070) );
  AOI22X1_RVT U3077 ( .A1(n1698), .A2(\read_value_mux[1][22] ), .A3(n1538), 
        .A4(\read_value_mux[1][23] ), .Y(n2043) );
  OA221X1_RVT U3078 ( .A1(n1538), .A2(\read_value_mux[1][23] ), .A3(n1699), 
        .A4(\read_value_mux[1][22] ), .A5(n2043), .Y(n2050) );
  AOI22X1_RVT U3079 ( .A1(n1701), .A2(\read_value_mux[1][20] ), .A3(n1703), 
        .A4(\read_value_mux[1][21] ), .Y(n2044) );
  OA221X1_RVT U3080 ( .A1(n1703), .A2(\read_value_mux[1][21] ), .A3(n1702), 
        .A4(\read_value_mux[1][20] ), .A5(n2044), .Y(n2049) );
  AOI22X1_RVT U3081 ( .A1(n1706), .A2(\read_value_mux[1][18] ), .A3(n1708), 
        .A4(\read_value_mux[1][19] ), .Y(n2045) );
  OA221X1_RVT U3082 ( .A1(n1708), .A2(\read_value_mux[1][19] ), .A3(n1706), 
        .A4(\read_value_mux[1][18] ), .A5(n2045), .Y(n2048) );
  AOI22X1_RVT U3083 ( .A1(n1710), .A2(\read_value_mux[1][16] ), .A3(n1713), 
        .A4(\read_value_mux[1][17] ), .Y(n2046) );
  OA221X1_RVT U3084 ( .A1(n1714), .A2(\read_value_mux[1][17] ), .A3(n1711), 
        .A4(\read_value_mux[1][16] ), .A5(n2046), .Y(n2047) );
  NAND4X0_RVT U3085 ( .A1(n2050), .A2(n2049), .A3(n2048), .A4(n2047), .Y(n2069) );
  AOI22X1_RVT U3086 ( .A1(n1716), .A2(\read_value_mux[1][14] ), .A3(n1718), 
        .A4(\read_value_mux[1][15] ), .Y(n2051) );
  OA221X1_RVT U3087 ( .A1(n1722), .A2(\read_value_mux[1][15] ), .A3(n1717), 
        .A4(\read_value_mux[1][14] ), .A5(n2051), .Y(n2058) );
  AOI22X1_RVT U3088 ( .A1(n1724), .A2(\read_value_mux[1][12] ), .A3(n1530), 
        .A4(\read_value_mux[1][13] ), .Y(n2052) );
  OA221X1_RVT U3089 ( .A1(n1530), .A2(\read_value_mux[1][13] ), .A3(n1725), 
        .A4(\read_value_mux[1][12] ), .A5(n2052), .Y(n2057) );
  AOI22X1_RVT U3090 ( .A1(n1728), .A2(\read_value_mux[1][10] ), .A3(n1730), 
        .A4(\read_value_mux[1][11] ), .Y(n2053) );
  OA221X1_RVT U3091 ( .A1(n1730), .A2(\read_value_mux[1][11] ), .A3(n1728), 
        .A4(\read_value_mux[1][10] ), .A5(n2053), .Y(n2056) );
  AOI22X1_RVT U3092 ( .A1(n1732), .A2(\read_value_mux[1][8] ), .A3(n1735), 
        .A4(\read_value_mux[1][9] ), .Y(n2054) );
  OA221X1_RVT U3093 ( .A1(n1736), .A2(\read_value_mux[1][9] ), .A3(n1733), 
        .A4(\read_value_mux[1][8] ), .A5(n2054), .Y(n2055) );
  NAND4X0_RVT U3094 ( .A1(n2058), .A2(n2057), .A3(n2056), .A4(n2055), .Y(n2068) );
  AOI22X1_RVT U3095 ( .A1(n1738), .A2(\read_value_mux[1][6] ), .A3(n1741), 
        .A4(\read_value_mux[1][7] ), .Y(n2059) );
  OA221X1_RVT U3096 ( .A1(n1740), .A2(\read_value_mux[1][7] ), .A3(n1738), 
        .A4(\read_value_mux[1][6] ), .A5(n2059), .Y(n2066) );
  AOI22X1_RVT U3097 ( .A1(n1742), .A2(\read_value_mux[1][4] ), .A3(n1744), 
        .A4(\read_value_mux[1][5] ), .Y(n2060) );
  OA221X1_RVT U3098 ( .A1(n1746), .A2(\read_value_mux[1][5] ), .A3(n1743), 
        .A4(\read_value_mux[1][4] ), .A5(n2060), .Y(n2065) );
  AOI22X1_RVT U3099 ( .A1(n1524), .A2(\read_value_mux[1][2] ), .A3(n1750), 
        .A4(\read_value_mux[1][3] ), .Y(n2061) );
  OA221X1_RVT U3100 ( .A1(n1750), .A2(\read_value_mux[1][3] ), .A3(n1748), 
        .A4(\read_value_mux[1][2] ), .A5(n2061), .Y(n2064) );
  OA221X1_RVT U3101 ( .A1(search_data[0]), .A2(n1667), .A3(n1752), .A4(
        \read_value_mux[1][0] ), .A5(search), .Y(n2062) );
  OA221X1_RVT U3102 ( .A1(search_data[31]), .A2(n1668), .A3(n1768), .A4(
        \read_value_mux[1][31] ), .A5(n2062), .Y(n2063) );
  NAND4X0_RVT U3103 ( .A1(n2066), .A2(n2065), .A3(n2064), .A4(n2063), .Y(n2067) );
  AO22X1_RVT U3104 ( .A1(search_data[28]), .A2(\read_value_mux[10][28] ), .A3(
        n1759), .A4(n1558), .Y(n2071) );
  OA221X1_RVT U3105 ( .A1(search_data[1]), .A2(n37), .A3(n1756), .A4(
        \read_value_mux[10][1] ), .A5(n2071), .Y(n2078) );
  AO22X1_RVT U3106 ( .A1(search_data[30]), .A2(\read_value_mux[10][30] ), .A3(
        n1765), .A4(n38), .Y(n2072) );
  OA221X1_RVT U3107 ( .A1(search_data[29]), .A2(n1669), .A3(n1762), .A4(
        \read_value_mux[10][29] ), .A5(n2072), .Y(n2077) );
  AOI22X1_RVT U3108 ( .A1(n1692), .A2(\read_value_mux[10][26] ), .A3(n1542), 
        .A4(\read_value_mux[10][27] ), .Y(n2073) );
  OA221X1_RVT U3109 ( .A1(n1542), .A2(\read_value_mux[10][27] ), .A3(n1691), 
        .A4(\read_value_mux[10][26] ), .A5(n2073), .Y(n2076) );
  AOI22X1_RVT U3110 ( .A1(n1696), .A2(\read_value_mux[10][24] ), .A3(n1540), 
        .A4(\read_value_mux[10][25] ), .Y(n2074) );
  OA221X1_RVT U3111 ( .A1(n1540), .A2(\read_value_mux[10][25] ), .A3(n1695), 
        .A4(\read_value_mux[10][24] ), .A5(n2074), .Y(n2075) );
  NAND4X0_RVT U3112 ( .A1(n2078), .A2(n2077), .A3(n2076), .A4(n2075), .Y(n2106) );
  AOI22X1_RVT U3113 ( .A1(n1699), .A2(\read_value_mux[10][22] ), .A3(n1538), 
        .A4(\read_value_mux[10][23] ), .Y(n2079) );
  OA221X1_RVT U3114 ( .A1(n1538), .A2(\read_value_mux[10][23] ), .A3(n1698), 
        .A4(\read_value_mux[10][22] ), .A5(n2079), .Y(n2086) );
  AOI22X1_RVT U3115 ( .A1(n1702), .A2(\read_value_mux[10][20] ), .A3(n1536), 
        .A4(\read_value_mux[10][21] ), .Y(n2080) );
  OA221X1_RVT U3116 ( .A1(n1703), .A2(\read_value_mux[10][21] ), .A3(n1701), 
        .A4(\read_value_mux[10][20] ), .A5(n2080), .Y(n2085) );
  AOI22X1_RVT U3117 ( .A1(n1706), .A2(\read_value_mux[10][18] ), .A3(n1534), 
        .A4(\read_value_mux[10][19] ), .Y(n2081) );
  OA221X1_RVT U3118 ( .A1(n1708), .A2(\read_value_mux[10][19] ), .A3(n1705), 
        .A4(\read_value_mux[10][18] ), .A5(n2081), .Y(n2084) );
  AOI22X1_RVT U3119 ( .A1(n1711), .A2(\read_value_mux[10][16] ), .A3(n1713), 
        .A4(\read_value_mux[10][17] ), .Y(n2082) );
  OA221X1_RVT U3120 ( .A1(n1714), .A2(\read_value_mux[10][17] ), .A3(n1710), 
        .A4(\read_value_mux[10][16] ), .A5(n2082), .Y(n2083) );
  NAND4X0_RVT U3121 ( .A1(n2086), .A2(n2085), .A3(n2084), .A4(n2083), .Y(n2105) );
  AOI22X1_RVT U3122 ( .A1(n1717), .A2(\read_value_mux[10][14] ), .A3(n1718), 
        .A4(\read_value_mux[10][15] ), .Y(n2087) );
  OA221X1_RVT U3123 ( .A1(n1722), .A2(\read_value_mux[10][15] ), .A3(n1716), 
        .A4(\read_value_mux[10][14] ), .A5(n2087), .Y(n2094) );
  AOI22X1_RVT U3124 ( .A1(n1725), .A2(\read_value_mux[10][12] ), .A3(n1530), 
        .A4(\read_value_mux[10][13] ), .Y(n2088) );
  OA221X1_RVT U3125 ( .A1(n1530), .A2(\read_value_mux[10][13] ), .A3(n1724), 
        .A4(\read_value_mux[10][12] ), .A5(n2088), .Y(n2093) );
  AOI22X1_RVT U3126 ( .A1(n1728), .A2(\read_value_mux[10][10] ), .A3(n1528), 
        .A4(\read_value_mux[10][11] ), .Y(n2089) );
  OA221X1_RVT U3127 ( .A1(n1730), .A2(\read_value_mux[10][11] ), .A3(n1727), 
        .A4(\read_value_mux[10][10] ), .A5(n2089), .Y(n2092) );
  AOI22X1_RVT U3128 ( .A1(n1733), .A2(\read_value_mux[10][8] ), .A3(n1735), 
        .A4(\read_value_mux[10][9] ), .Y(n2090) );
  OA221X1_RVT U3129 ( .A1(n1736), .A2(\read_value_mux[10][9] ), .A3(n1732), 
        .A4(\read_value_mux[10][8] ), .A5(n2090), .Y(n2091) );
  NAND4X0_RVT U3130 ( .A1(n2094), .A2(n2093), .A3(n2092), .A4(n2091), .Y(n2104) );
  AOI22X1_RVT U3131 ( .A1(n1738), .A2(\read_value_mux[10][6] ), .A3(n1740), 
        .A4(\read_value_mux[10][7] ), .Y(n2095) );
  OA221X1_RVT U3132 ( .A1(n1740), .A2(\read_value_mux[10][7] ), .A3(n1738), 
        .A4(\read_value_mux[10][6] ), .A5(n2095), .Y(n2102) );
  AOI22X1_RVT U3133 ( .A1(n1743), .A2(\read_value_mux[10][4] ), .A3(n1744), 
        .A4(\read_value_mux[10][5] ), .Y(n2096) );
  OA221X1_RVT U3134 ( .A1(n1746), .A2(\read_value_mux[10][5] ), .A3(n1742), 
        .A4(\read_value_mux[10][4] ), .A5(n2096), .Y(n2101) );
  AOI22X1_RVT U3135 ( .A1(n1748), .A2(\read_value_mux[10][2] ), .A3(n1750), 
        .A4(\read_value_mux[10][3] ), .Y(n2097) );
  OA221X1_RVT U3136 ( .A1(n1750), .A2(\read_value_mux[10][3] ), .A3(n1524), 
        .A4(\read_value_mux[10][2] ), .A5(n2097), .Y(n2100) );
  OA221X1_RVT U3137 ( .A1(search_data[0]), .A2(n1602), .A3(n1753), .A4(
        \read_value_mux[10][0] ), .A5(search), .Y(n2098) );
  OA221X1_RVT U3138 ( .A1(search_data[31]), .A2(n1670), .A3(n1768), .A4(
        \read_value_mux[10][31] ), .A5(n2098), .Y(n2099) );
  NAND4X0_RVT U3139 ( .A1(n2102), .A2(n2101), .A3(n2100), .A4(n2099), .Y(n2103) );
  AO22X1_RVT U3140 ( .A1(search_data[28]), .A2(\read_value_mux[12][28] ), .A3(
        n1758), .A4(n1545), .Y(n2107) );
  OA221X1_RVT U3141 ( .A1(search_data[1]), .A2(n43), .A3(n1755), .A4(
        \read_value_mux[12][1] ), .A5(n2107), .Y(n2114) );
  AO22X1_RVT U3142 ( .A1(search_data[30]), .A2(\read_value_mux[12][30] ), .A3(
        n1764), .A4(n44), .Y(n2108) );
  OA221X1_RVT U3143 ( .A1(search_data[29]), .A2(n1569), .A3(n1762), .A4(
        \read_value_mux[12][29] ), .A5(n2108), .Y(n2113) );
  AOI22X1_RVT U3144 ( .A1(n1543), .A2(\read_value_mux[12][26] ), .A3(n1542), 
        .A4(\read_value_mux[12][27] ), .Y(n2109) );
  OA221X1_RVT U3145 ( .A1(n1542), .A2(\read_value_mux[12][27] ), .A3(n1692), 
        .A4(\read_value_mux[12][26] ), .A5(n2109), .Y(n2112) );
  AOI22X1_RVT U3146 ( .A1(n1541), .A2(\read_value_mux[12][24] ), .A3(n1540), 
        .A4(\read_value_mux[12][25] ), .Y(n2110) );
  OA221X1_RVT U3147 ( .A1(n1540), .A2(\read_value_mux[12][25] ), .A3(n1696), 
        .A4(\read_value_mux[12][24] ), .A5(n2110), .Y(n2111) );
  NAND4X0_RVT U3148 ( .A1(n2114), .A2(n2113), .A3(n2112), .A4(n2111), .Y(n2142) );
  AOI22X1_RVT U3149 ( .A1(n1539), .A2(\read_value_mux[12][22] ), .A3(n1538), 
        .A4(\read_value_mux[12][23] ), .Y(n2115) );
  OA221X1_RVT U3150 ( .A1(n1538), .A2(\read_value_mux[12][23] ), .A3(n1699), 
        .A4(\read_value_mux[12][22] ), .A5(n2115), .Y(n2122) );
  AOI22X1_RVT U3151 ( .A1(n1537), .A2(\read_value_mux[12][20] ), .A3(n1536), 
        .A4(\read_value_mux[12][21] ), .Y(n2116) );
  OA221X1_RVT U3152 ( .A1(n1536), .A2(\read_value_mux[12][21] ), .A3(n1702), 
        .A4(\read_value_mux[12][20] ), .A5(n2116), .Y(n2121) );
  AOI22X1_RVT U3153 ( .A1(n1535), .A2(\read_value_mux[12][18] ), .A3(n1534), 
        .A4(\read_value_mux[12][19] ), .Y(n2117) );
  OA221X1_RVT U3154 ( .A1(n1534), .A2(\read_value_mux[12][19] ), .A3(n1706), 
        .A4(\read_value_mux[12][18] ), .A5(n2117), .Y(n2120) );
  AOI22X1_RVT U3155 ( .A1(n1533), .A2(\read_value_mux[12][16] ), .A3(n1713), 
        .A4(\read_value_mux[12][17] ), .Y(n2118) );
  OA221X1_RVT U3156 ( .A1(n1713), .A2(\read_value_mux[12][17] ), .A3(n1711), 
        .A4(\read_value_mux[12][16] ), .A5(n2118), .Y(n2119) );
  NAND4X0_RVT U3157 ( .A1(n2122), .A2(n2121), .A3(n2120), .A4(n2119), .Y(n2141) );
  AOI22X1_RVT U3158 ( .A1(n1532), .A2(\read_value_mux[12][14] ), .A3(n1718), 
        .A4(\read_value_mux[12][15] ), .Y(n2123) );
  OA221X1_RVT U3159 ( .A1(n1721), .A2(\read_value_mux[12][15] ), .A3(n1717), 
        .A4(\read_value_mux[12][14] ), .A5(n2123), .Y(n2130) );
  AOI22X1_RVT U3160 ( .A1(n1531), .A2(\read_value_mux[12][12] ), .A3(n1530), 
        .A4(\read_value_mux[12][13] ), .Y(n2124) );
  OA221X1_RVT U3161 ( .A1(n1530), .A2(\read_value_mux[12][13] ), .A3(n1725), 
        .A4(\read_value_mux[12][12] ), .A5(n2124), .Y(n2129) );
  AOI22X1_RVT U3162 ( .A1(n1529), .A2(\read_value_mux[12][10] ), .A3(n1528), 
        .A4(\read_value_mux[12][11] ), .Y(n2125) );
  OA221X1_RVT U3163 ( .A1(n1528), .A2(\read_value_mux[12][11] ), .A3(n1728), 
        .A4(\read_value_mux[12][10] ), .A5(n2125), .Y(n2128) );
  AOI22X1_RVT U3164 ( .A1(n1527), .A2(\read_value_mux[12][8] ), .A3(n1735), 
        .A4(\read_value_mux[12][9] ), .Y(n2126) );
  OA221X1_RVT U3165 ( .A1(n1735), .A2(\read_value_mux[12][9] ), .A3(n1733), 
        .A4(\read_value_mux[12][8] ), .A5(n2126), .Y(n2127) );
  NAND4X0_RVT U3166 ( .A1(n2130), .A2(n2129), .A3(n2128), .A4(n2127), .Y(n2140) );
  AOI22X1_RVT U3167 ( .A1(n2940), .A2(\read_value_mux[12][6] ), .A3(n1739), 
        .A4(\read_value_mux[12][7] ), .Y(n2131) );
  OA221X1_RVT U3168 ( .A1(n1740), .A2(\read_value_mux[12][7] ), .A3(n1738), 
        .A4(\read_value_mux[12][6] ), .A5(n2131), .Y(n2138) );
  AOI22X1_RVT U3169 ( .A1(n1526), .A2(\read_value_mux[12][4] ), .A3(n1744), 
        .A4(\read_value_mux[12][5] ), .Y(n2132) );
  OA221X1_RVT U3170 ( .A1(n1745), .A2(\read_value_mux[12][5] ), .A3(n1743), 
        .A4(\read_value_mux[12][4] ), .A5(n2132), .Y(n2137) );
  AOI22X1_RVT U3171 ( .A1(n1524), .A2(\read_value_mux[12][2] ), .A3(n1750), 
        .A4(\read_value_mux[12][3] ), .Y(n2133) );
  OA221X1_RVT U3172 ( .A1(n1750), .A2(\read_value_mux[12][3] ), .A3(n1748), 
        .A4(\read_value_mux[12][2] ), .A5(n2133), .Y(n2136) );
  OA221X1_RVT U3173 ( .A1(search_data[0]), .A2(n1570), .A3(n1752), .A4(
        \read_value_mux[12][0] ), .A5(search), .Y(n2134) );
  OA221X1_RVT U3174 ( .A1(search_data[31]), .A2(n1571), .A3(n1768), .A4(
        \read_value_mux[12][31] ), .A5(n2134), .Y(n2135) );
  NAND4X0_RVT U3175 ( .A1(n2138), .A2(n2137), .A3(n2136), .A4(n2135), .Y(n2139) );
  AO22X1_RVT U3176 ( .A1(search_data[28]), .A2(\read_value_mux[13][28] ), .A3(
        n1758), .A4(n1559), .Y(n2143) );
  OA221X1_RVT U3177 ( .A1(search_data[1]), .A2(n45), .A3(n1755), .A4(
        \read_value_mux[13][1] ), .A5(n2143), .Y(n2150) );
  AO22X1_RVT U3178 ( .A1(search_data[30]), .A2(\read_value_mux[13][30] ), .A3(
        n1764), .A4(n46), .Y(n2144) );
  OA221X1_RVT U3179 ( .A1(search_data[29]), .A2(n1603), .A3(n1761), .A4(
        \read_value_mux[13][29] ), .A5(n2144), .Y(n2149) );
  AOI22X1_RVT U3180 ( .A1(n1543), .A2(\read_value_mux[13][26] ), .A3(n1542), 
        .A4(\read_value_mux[13][27] ), .Y(n2145) );
  OA221X1_RVT U3181 ( .A1(n1542), .A2(\read_value_mux[13][27] ), .A3(n1691), 
        .A4(\read_value_mux[13][26] ), .A5(n2145), .Y(n2148) );
  AOI22X1_RVT U3182 ( .A1(n1541), .A2(\read_value_mux[13][24] ), .A3(n1697), 
        .A4(\read_value_mux[13][25] ), .Y(n2146) );
  OA221X1_RVT U3183 ( .A1(n1540), .A2(\read_value_mux[13][25] ), .A3(n1695), 
        .A4(\read_value_mux[13][24] ), .A5(n2146), .Y(n2147) );
  NAND4X0_RVT U3184 ( .A1(n2150), .A2(n2149), .A3(n2148), .A4(n2147), .Y(n2178) );
  AOI22X1_RVT U3185 ( .A1(n1539), .A2(\read_value_mux[13][22] ), .A3(n1538), 
        .A4(\read_value_mux[13][23] ), .Y(n2151) );
  OA221X1_RVT U3186 ( .A1(n1538), .A2(\read_value_mux[13][23] ), .A3(n1698), 
        .A4(\read_value_mux[13][22] ), .A5(n2151), .Y(n2158) );
  AOI22X1_RVT U3187 ( .A1(n1537), .A2(\read_value_mux[13][20] ), .A3(n1536), 
        .A4(\read_value_mux[13][21] ), .Y(n2152) );
  OA221X1_RVT U3188 ( .A1(n1703), .A2(\read_value_mux[13][21] ), .A3(n1701), 
        .A4(\read_value_mux[13][20] ), .A5(n2152), .Y(n2157) );
  AOI22X1_RVT U3189 ( .A1(n1535), .A2(\read_value_mux[13][18] ), .A3(n1534), 
        .A4(\read_value_mux[13][19] ), .Y(n2153) );
  OA221X1_RVT U3190 ( .A1(n1708), .A2(\read_value_mux[13][19] ), .A3(n1705), 
        .A4(\read_value_mux[13][18] ), .A5(n2153), .Y(n2156) );
  AOI22X1_RVT U3191 ( .A1(n1533), .A2(\read_value_mux[13][16] ), .A3(n1713), 
        .A4(\read_value_mux[13][17] ), .Y(n2154) );
  OA221X1_RVT U3192 ( .A1(n1714), .A2(\read_value_mux[13][17] ), .A3(n1710), 
        .A4(\read_value_mux[13][16] ), .A5(n2154), .Y(n2155) );
  NAND4X0_RVT U3193 ( .A1(n2158), .A2(n2157), .A3(n2156), .A4(n2155), .Y(n2177) );
  AOI22X1_RVT U3194 ( .A1(n1532), .A2(\read_value_mux[13][14] ), .A3(n1718), 
        .A4(\read_value_mux[13][15] ), .Y(n2159) );
  OA221X1_RVT U3195 ( .A1(n1722), .A2(\read_value_mux[13][15] ), .A3(n1716), 
        .A4(\read_value_mux[13][14] ), .A5(n2159), .Y(n2166) );
  AOI22X1_RVT U3196 ( .A1(n1531), .A2(\read_value_mux[13][12] ), .A3(n1530), 
        .A4(\read_value_mux[13][13] ), .Y(n2160) );
  OA221X1_RVT U3197 ( .A1(n1530), .A2(\read_value_mux[13][13] ), .A3(n1724), 
        .A4(\read_value_mux[13][12] ), .A5(n2160), .Y(n2165) );
  AOI22X1_RVT U3198 ( .A1(n1529), .A2(\read_value_mux[13][10] ), .A3(n1528), 
        .A4(\read_value_mux[13][11] ), .Y(n2161) );
  OA221X1_RVT U3199 ( .A1(n1730), .A2(\read_value_mux[13][11] ), .A3(n1727), 
        .A4(\read_value_mux[13][10] ), .A5(n2161), .Y(n2164) );
  AOI22X1_RVT U3200 ( .A1(n1527), .A2(\read_value_mux[13][8] ), .A3(n1735), 
        .A4(\read_value_mux[13][9] ), .Y(n2162) );
  OA221X1_RVT U3201 ( .A1(n1736), .A2(\read_value_mux[13][9] ), .A3(n1732), 
        .A4(\read_value_mux[13][8] ), .A5(n2162), .Y(n2163) );
  NAND4X0_RVT U3202 ( .A1(n2166), .A2(n2165), .A3(n2164), .A4(n2163), .Y(n2176) );
  AOI22X1_RVT U3203 ( .A1(n2940), .A2(\read_value_mux[13][6] ), .A3(n1741), 
        .A4(\read_value_mux[13][7] ), .Y(n2167) );
  OA221X1_RVT U3204 ( .A1(n1740), .A2(\read_value_mux[13][7] ), .A3(n1738), 
        .A4(\read_value_mux[13][6] ), .A5(n2167), .Y(n2174) );
  AOI22X1_RVT U3205 ( .A1(n1526), .A2(\read_value_mux[13][4] ), .A3(n1744), 
        .A4(\read_value_mux[13][5] ), .Y(n2168) );
  OA221X1_RVT U3206 ( .A1(n1746), .A2(\read_value_mux[13][5] ), .A3(n1742), 
        .A4(\read_value_mux[13][4] ), .A5(n2168), .Y(n2173) );
  AOI22X1_RVT U3207 ( .A1(n1524), .A2(\read_value_mux[13][2] ), .A3(n1750), 
        .A4(\read_value_mux[13][3] ), .Y(n2169) );
  OA221X1_RVT U3208 ( .A1(n1750), .A2(\read_value_mux[13][3] ), .A3(n1524), 
        .A4(\read_value_mux[13][2] ), .A5(n2169), .Y(n2172) );
  OA221X1_RVT U3209 ( .A1(search_data[0]), .A2(n1604), .A3(n1752), .A4(
        \read_value_mux[13][0] ), .A5(search), .Y(n2170) );
  OA221X1_RVT U3210 ( .A1(search_data[31]), .A2(n1605), .A3(n1767), .A4(
        \read_value_mux[13][31] ), .A5(n2170), .Y(n2171) );
  NAND4X0_RVT U3211 ( .A1(n2174), .A2(n2173), .A3(n2172), .A4(n2171), .Y(n2175) );
  AO22X1_RVT U3212 ( .A1(search_data[28]), .A2(\read_value_mux[16][28] ), .A3(
        n1758), .A4(n1546), .Y(n2179) );
  OA221X1_RVT U3213 ( .A1(search_data[1]), .A2(n53), .A3(n1755), .A4(
        \read_value_mux[16][1] ), .A5(n2179), .Y(n2186) );
  AO22X1_RVT U3214 ( .A1(search_data[30]), .A2(\read_value_mux[16][30] ), .A3(
        n1764), .A4(n54), .Y(n2180) );
  OA221X1_RVT U3215 ( .A1(search_data[29]), .A2(n1572), .A3(n1761), .A4(
        \read_value_mux[16][29] ), .A5(n2180), .Y(n2185) );
  AOI22X1_RVT U3216 ( .A1(n1543), .A2(\read_value_mux[16][26] ), .A3(n1694), 
        .A4(\read_value_mux[16][27] ), .Y(n2181) );
  OA221X1_RVT U3217 ( .A1(n1542), .A2(\read_value_mux[16][27] ), .A3(n1691), 
        .A4(\read_value_mux[16][26] ), .A5(n2181), .Y(n2184) );
  AOI22X1_RVT U3218 ( .A1(n1541), .A2(\read_value_mux[16][24] ), .A3(n1697), 
        .A4(\read_value_mux[16][25] ), .Y(n2182) );
  OA221X1_RVT U3219 ( .A1(n1540), .A2(\read_value_mux[16][25] ), .A3(n1695), 
        .A4(\read_value_mux[16][24] ), .A5(n2182), .Y(n2183) );
  NAND4X0_RVT U3220 ( .A1(n2186), .A2(n2185), .A3(n2184), .A4(n2183), .Y(n2214) );
  AOI22X1_RVT U3221 ( .A1(n1539), .A2(\read_value_mux[16][22] ), .A3(n1700), 
        .A4(\read_value_mux[16][23] ), .Y(n2187) );
  OA221X1_RVT U3222 ( .A1(n1538), .A2(\read_value_mux[16][23] ), .A3(n1698), 
        .A4(\read_value_mux[16][22] ), .A5(n2187), .Y(n2194) );
  AOI22X1_RVT U3223 ( .A1(n1537), .A2(\read_value_mux[16][20] ), .A3(n1536), 
        .A4(\read_value_mux[16][21] ), .Y(n2188) );
  OA221X1_RVT U3224 ( .A1(n1536), .A2(\read_value_mux[16][21] ), .A3(n1701), 
        .A4(\read_value_mux[16][20] ), .A5(n2188), .Y(n2193) );
  AOI22X1_RVT U3225 ( .A1(n1535), .A2(\read_value_mux[16][18] ), .A3(n1534), 
        .A4(\read_value_mux[16][19] ), .Y(n2189) );
  OA221X1_RVT U3226 ( .A1(n1534), .A2(\read_value_mux[16][19] ), .A3(n1705), 
        .A4(\read_value_mux[16][18] ), .A5(n2189), .Y(n2192) );
  AOI22X1_RVT U3227 ( .A1(n1533), .A2(\read_value_mux[16][16] ), .A3(n1712), 
        .A4(\read_value_mux[16][17] ), .Y(n2190) );
  OA221X1_RVT U3228 ( .A1(n1713), .A2(\read_value_mux[16][17] ), .A3(n1710), 
        .A4(\read_value_mux[16][16] ), .A5(n2190), .Y(n2191) );
  NAND4X0_RVT U3229 ( .A1(n2194), .A2(n2193), .A3(n2192), .A4(n2191), .Y(n2213) );
  AOI22X1_RVT U3230 ( .A1(n1532), .A2(\read_value_mux[16][14] ), .A3(n1718), 
        .A4(\read_value_mux[16][15] ), .Y(n2195) );
  OA221X1_RVT U3231 ( .A1(n1721), .A2(\read_value_mux[16][15] ), .A3(n1716), 
        .A4(\read_value_mux[16][14] ), .A5(n2195), .Y(n2202) );
  AOI22X1_RVT U3232 ( .A1(n1531), .A2(\read_value_mux[16][12] ), .A3(n1726), 
        .A4(\read_value_mux[16][13] ), .Y(n2196) );
  OA221X1_RVT U3233 ( .A1(n1530), .A2(\read_value_mux[16][13] ), .A3(n1724), 
        .A4(\read_value_mux[16][12] ), .A5(n2196), .Y(n2201) );
  AOI22X1_RVT U3234 ( .A1(n1529), .A2(\read_value_mux[16][10] ), .A3(n1528), 
        .A4(\read_value_mux[16][11] ), .Y(n2197) );
  OA221X1_RVT U3235 ( .A1(n1528), .A2(\read_value_mux[16][11] ), .A3(n1727), 
        .A4(\read_value_mux[16][10] ), .A5(n2197), .Y(n2200) );
  AOI22X1_RVT U3236 ( .A1(n1527), .A2(\read_value_mux[16][8] ), .A3(n1734), 
        .A4(\read_value_mux[16][9] ), .Y(n2198) );
  OA221X1_RVT U3237 ( .A1(n1735), .A2(\read_value_mux[16][9] ), .A3(n1732), 
        .A4(\read_value_mux[16][8] ), .A5(n2198), .Y(n2199) );
  NAND4X0_RVT U3238 ( .A1(n2202), .A2(n2201), .A3(n2200), .A4(n2199), .Y(n2212) );
  AOI22X1_RVT U3239 ( .A1(n2940), .A2(\read_value_mux[16][6] ), .A3(n1741), 
        .A4(\read_value_mux[16][7] ), .Y(n2203) );
  OA221X1_RVT U3240 ( .A1(n1740), .A2(\read_value_mux[16][7] ), .A3(n1738), 
        .A4(\read_value_mux[16][6] ), .A5(n2203), .Y(n2210) );
  AOI22X1_RVT U3241 ( .A1(n1526), .A2(\read_value_mux[16][4] ), .A3(n1744), 
        .A4(\read_value_mux[16][5] ), .Y(n2204) );
  OA221X1_RVT U3242 ( .A1(n1745), .A2(\read_value_mux[16][5] ), .A3(n1742), 
        .A4(\read_value_mux[16][4] ), .A5(n2204), .Y(n2209) );
  AOI22X1_RVT U3243 ( .A1(n1524), .A2(\read_value_mux[16][2] ), .A3(n1750), 
        .A4(\read_value_mux[16][3] ), .Y(n2205) );
  OA221X1_RVT U3244 ( .A1(n1750), .A2(\read_value_mux[16][3] ), .A3(n1524), 
        .A4(\read_value_mux[16][2] ), .A5(n2205), .Y(n2208) );
  OA221X1_RVT U3245 ( .A1(search_data[0]), .A2(n1573), .A3(n1752), .A4(
        \read_value_mux[16][0] ), .A5(search), .Y(n2206) );
  OA221X1_RVT U3246 ( .A1(search_data[31]), .A2(n1574), .A3(n1767), .A4(
        \read_value_mux[16][31] ), .A5(n2206), .Y(n2207) );
  NAND4X0_RVT U3247 ( .A1(n2210), .A2(n2209), .A3(n2208), .A4(n2207), .Y(n2211) );
  AO22X1_RVT U3248 ( .A1(search_data[28]), .A2(\read_value_mux[18][28] ), .A3(
        n1758), .A4(n1560), .Y(n2215) );
  OA221X1_RVT U3249 ( .A1(search_data[1]), .A2(n58), .A3(n1755), .A4(
        \read_value_mux[18][1] ), .A5(n2215), .Y(n2222) );
  AO22X1_RVT U3250 ( .A1(search_data[30]), .A2(\read_value_mux[18][30] ), .A3(
        n1764), .A4(n59), .Y(n2216) );
  OA221X1_RVT U3251 ( .A1(search_data[29]), .A2(n1606), .A3(n1761), .A4(
        \read_value_mux[18][29] ), .A5(n2216), .Y(n2221) );
  AOI22X1_RVT U3252 ( .A1(n1543), .A2(\read_value_mux[18][26] ), .A3(n1694), 
        .A4(\read_value_mux[18][27] ), .Y(n2217) );
  OA221X1_RVT U3253 ( .A1(n1542), .A2(\read_value_mux[18][27] ), .A3(n1692), 
        .A4(\read_value_mux[18][26] ), .A5(n2217), .Y(n2220) );
  AOI22X1_RVT U3254 ( .A1(n1541), .A2(\read_value_mux[18][24] ), .A3(n1540), 
        .A4(\read_value_mux[18][25] ), .Y(n2218) );
  OA221X1_RVT U3255 ( .A1(n1540), .A2(\read_value_mux[18][25] ), .A3(n1696), 
        .A4(\read_value_mux[18][24] ), .A5(n2218), .Y(n2219) );
  NAND4X0_RVT U3256 ( .A1(n2222), .A2(n2221), .A3(n2220), .A4(n2219), .Y(n2250) );
  AOI22X1_RVT U3257 ( .A1(n1539), .A2(\read_value_mux[18][22] ), .A3(n1700), 
        .A4(\read_value_mux[18][23] ), .Y(n2223) );
  OA221X1_RVT U3258 ( .A1(n1538), .A2(\read_value_mux[18][23] ), .A3(n1699), 
        .A4(\read_value_mux[18][22] ), .A5(n2223), .Y(n2230) );
  AOI22X1_RVT U3259 ( .A1(n1537), .A2(\read_value_mux[18][20] ), .A3(n1536), 
        .A4(\read_value_mux[18][21] ), .Y(n2224) );
  OA221X1_RVT U3260 ( .A1(n1703), .A2(\read_value_mux[18][21] ), .A3(n1702), 
        .A4(\read_value_mux[18][20] ), .A5(n2224), .Y(n2229) );
  AOI22X1_RVT U3261 ( .A1(n1535), .A2(\read_value_mux[18][18] ), .A3(n1534), 
        .A4(\read_value_mux[18][19] ), .Y(n2225) );
  OA221X1_RVT U3262 ( .A1(n1708), .A2(\read_value_mux[18][19] ), .A3(n1706), 
        .A4(\read_value_mux[18][18] ), .A5(n2225), .Y(n2228) );
  AOI22X1_RVT U3263 ( .A1(n1533), .A2(\read_value_mux[18][16] ), .A3(n1713), 
        .A4(\read_value_mux[18][17] ), .Y(n2226) );
  OA221X1_RVT U3264 ( .A1(n1714), .A2(\read_value_mux[18][17] ), .A3(n1711), 
        .A4(\read_value_mux[18][16] ), .A5(n2226), .Y(n2227) );
  NAND4X0_RVT U3265 ( .A1(n2230), .A2(n2229), .A3(n2228), .A4(n2227), .Y(n2249) );
  AOI22X1_RVT U3266 ( .A1(n1532), .A2(\read_value_mux[18][14] ), .A3(n1718), 
        .A4(\read_value_mux[18][15] ), .Y(n2231) );
  OA221X1_RVT U3267 ( .A1(n1721), .A2(\read_value_mux[18][15] ), .A3(n1717), 
        .A4(\read_value_mux[18][14] ), .A5(n2231), .Y(n2238) );
  AOI22X1_RVT U3268 ( .A1(n1531), .A2(\read_value_mux[18][12] ), .A3(n1726), 
        .A4(\read_value_mux[18][13] ), .Y(n2232) );
  OA221X1_RVT U3269 ( .A1(n1530), .A2(\read_value_mux[18][13] ), .A3(n1725), 
        .A4(\read_value_mux[18][12] ), .A5(n2232), .Y(n2237) );
  AOI22X1_RVT U3270 ( .A1(n1529), .A2(\read_value_mux[18][10] ), .A3(n1528), 
        .A4(\read_value_mux[18][11] ), .Y(n2233) );
  OA221X1_RVT U3271 ( .A1(n1730), .A2(\read_value_mux[18][11] ), .A3(n1728), 
        .A4(\read_value_mux[18][10] ), .A5(n2233), .Y(n2236) );
  AOI22X1_RVT U3272 ( .A1(n1527), .A2(\read_value_mux[18][8] ), .A3(n1735), 
        .A4(\read_value_mux[18][9] ), .Y(n2234) );
  OA221X1_RVT U3273 ( .A1(n1736), .A2(\read_value_mux[18][9] ), .A3(n1733), 
        .A4(\read_value_mux[18][8] ), .A5(n2234), .Y(n2235) );
  NAND4X0_RVT U3274 ( .A1(n2238), .A2(n2237), .A3(n2236), .A4(n2235), .Y(n2248) );
  AOI22X1_RVT U3275 ( .A1(n2940), .A2(\read_value_mux[18][6] ), .A3(n1741), 
        .A4(\read_value_mux[18][7] ), .Y(n2239) );
  OA221X1_RVT U3276 ( .A1(n1740), .A2(\read_value_mux[18][7] ), .A3(n1738), 
        .A4(\read_value_mux[18][6] ), .A5(n2239), .Y(n2246) );
  AOI22X1_RVT U3277 ( .A1(n1526), .A2(\read_value_mux[18][4] ), .A3(n1744), 
        .A4(\read_value_mux[18][5] ), .Y(n2240) );
  OA221X1_RVT U3278 ( .A1(n1745), .A2(\read_value_mux[18][5] ), .A3(n1743), 
        .A4(\read_value_mux[18][4] ), .A5(n2240), .Y(n2245) );
  AOI22X1_RVT U3279 ( .A1(n1524), .A2(\read_value_mux[18][2] ), .A3(n1750), 
        .A4(\read_value_mux[18][3] ), .Y(n2241) );
  OA221X1_RVT U3280 ( .A1(n1750), .A2(\read_value_mux[18][3] ), .A3(n1748), 
        .A4(\read_value_mux[18][2] ), .A5(n2241), .Y(n2244) );
  OA221X1_RVT U3281 ( .A1(search_data[0]), .A2(n1607), .A3(n1752), .A4(
        \read_value_mux[18][0] ), .A5(search), .Y(n2242) );
  OA221X1_RVT U3282 ( .A1(search_data[31]), .A2(n1608), .A3(n1767), .A4(
        \read_value_mux[18][31] ), .A5(n2242), .Y(n2243) );
  NAND4X0_RVT U3283 ( .A1(n2246), .A2(n2245), .A3(n2244), .A4(n2243), .Y(n2247) );
  OR4X1_RVT U3284 ( .A1(n2250), .A2(n2249), .A3(n2248), .A4(n2247), .Y(n2983)
         );
  NAND2X0_RVT U3285 ( .A1(n2985), .A2(n2983), .Y(n2653) );
  AO22X1_RVT U3286 ( .A1(search_data[28]), .A2(\read_value_mux[19][28] ), .A3(
        n1758), .A4(n1547), .Y(n2251) );
  OA221X1_RVT U3287 ( .A1(search_data[1]), .A2(n60), .A3(n1755), .A4(
        \read_value_mux[19][1] ), .A5(n2251), .Y(n2258) );
  AO22X1_RVT U3288 ( .A1(search_data[30]), .A2(\read_value_mux[19][30] ), .A3(
        n1764), .A4(n61), .Y(n2252) );
  OA221X1_RVT U3289 ( .A1(search_data[29]), .A2(n1654), .A3(n1761), .A4(
        \read_value_mux[19][29] ), .A5(n2252), .Y(n2257) );
  AOI22X1_RVT U3290 ( .A1(n1543), .A2(\read_value_mux[19][26] ), .A3(n1542), 
        .A4(\read_value_mux[19][27] ), .Y(n2253) );
  OA221X1_RVT U3291 ( .A1(n1542), .A2(\read_value_mux[19][27] ), .A3(n1691), 
        .A4(\read_value_mux[19][26] ), .A5(n2253), .Y(n2256) );
  AOI22X1_RVT U3292 ( .A1(n1541), .A2(\read_value_mux[19][24] ), .A3(n1540), 
        .A4(\read_value_mux[19][25] ), .Y(n2254) );
  OA221X1_RVT U3293 ( .A1(n1540), .A2(\read_value_mux[19][25] ), .A3(n1696), 
        .A4(\read_value_mux[19][24] ), .A5(n2254), .Y(n2255) );
  NAND4X0_RVT U3294 ( .A1(n2258), .A2(n2257), .A3(n2256), .A4(n2255), .Y(n2286) );
  AOI22X1_RVT U3295 ( .A1(n1539), .A2(\read_value_mux[19][22] ), .A3(n1538), 
        .A4(\read_value_mux[19][23] ), .Y(n2259) );
  OA221X1_RVT U3296 ( .A1(n1538), .A2(\read_value_mux[19][23] ), .A3(n1699), 
        .A4(\read_value_mux[19][22] ), .A5(n2259), .Y(n2266) );
  AOI22X1_RVT U3297 ( .A1(n1537), .A2(\read_value_mux[19][20] ), .A3(n1536), 
        .A4(\read_value_mux[19][21] ), .Y(n2260) );
  OA221X1_RVT U3298 ( .A1(n1703), .A2(\read_value_mux[19][21] ), .A3(n1702), 
        .A4(\read_value_mux[19][20] ), .A5(n2260), .Y(n2265) );
  AOI22X1_RVT U3299 ( .A1(n1535), .A2(\read_value_mux[19][18] ), .A3(n1534), 
        .A4(\read_value_mux[19][19] ), .Y(n2261) );
  OA221X1_RVT U3300 ( .A1(n1708), .A2(\read_value_mux[19][19] ), .A3(n1705), 
        .A4(\read_value_mux[19][18] ), .A5(n2261), .Y(n2264) );
  AOI22X1_RVT U3301 ( .A1(n1533), .A2(\read_value_mux[19][16] ), .A3(n1712), 
        .A4(\read_value_mux[19][17] ), .Y(n2262) );
  OA221X1_RVT U3302 ( .A1(n1714), .A2(\read_value_mux[19][17] ), .A3(n1711), 
        .A4(\read_value_mux[19][16] ), .A5(n2262), .Y(n2263) );
  NAND4X0_RVT U3303 ( .A1(n2266), .A2(n2265), .A3(n2264), .A4(n2263), .Y(n2285) );
  AOI22X1_RVT U3304 ( .A1(n1532), .A2(\read_value_mux[19][14] ), .A3(n1719), 
        .A4(\read_value_mux[19][15] ), .Y(n2267) );
  OA221X1_RVT U3305 ( .A1(n1721), .A2(\read_value_mux[19][15] ), .A3(n1717), 
        .A4(\read_value_mux[19][14] ), .A5(n2267), .Y(n2274) );
  AOI22X1_RVT U3306 ( .A1(n1531), .A2(\read_value_mux[19][12] ), .A3(n1530), 
        .A4(\read_value_mux[19][13] ), .Y(n2268) );
  OA221X1_RVT U3307 ( .A1(n1530), .A2(\read_value_mux[19][13] ), .A3(n1725), 
        .A4(\read_value_mux[19][12] ), .A5(n2268), .Y(n2273) );
  AOI22X1_RVT U3308 ( .A1(n1529), .A2(\read_value_mux[19][10] ), .A3(n1528), 
        .A4(\read_value_mux[19][11] ), .Y(n2269) );
  OA221X1_RVT U3309 ( .A1(n1730), .A2(\read_value_mux[19][11] ), .A3(n1727), 
        .A4(\read_value_mux[19][10] ), .A5(n2269), .Y(n2272) );
  AOI22X1_RVT U3310 ( .A1(n1527), .A2(\read_value_mux[19][8] ), .A3(n1734), 
        .A4(\read_value_mux[19][9] ), .Y(n2270) );
  OA221X1_RVT U3311 ( .A1(n1736), .A2(\read_value_mux[19][9] ), .A3(n1733), 
        .A4(\read_value_mux[19][8] ), .A5(n2270), .Y(n2271) );
  NAND4X0_RVT U3312 ( .A1(n2274), .A2(n2273), .A3(n2272), .A4(n2271), .Y(n2284) );
  AOI22X1_RVT U3313 ( .A1(n2940), .A2(\read_value_mux[19][6] ), .A3(n1741), 
        .A4(\read_value_mux[19][7] ), .Y(n2275) );
  OA221X1_RVT U3314 ( .A1(n1740), .A2(\read_value_mux[19][7] ), .A3(n1738), 
        .A4(\read_value_mux[19][6] ), .A5(n2275), .Y(n2282) );
  AOI22X1_RVT U3315 ( .A1(n1526), .A2(\read_value_mux[19][4] ), .A3(n1525), 
        .A4(\read_value_mux[19][5] ), .Y(n2276) );
  OA221X1_RVT U3316 ( .A1(n1745), .A2(\read_value_mux[19][5] ), .A3(n1743), 
        .A4(\read_value_mux[19][4] ), .A5(n2276), .Y(n2281) );
  AOI22X1_RVT U3317 ( .A1(n1524), .A2(\read_value_mux[19][2] ), .A3(n1750), 
        .A4(\read_value_mux[19][3] ), .Y(n2277) );
  OA221X1_RVT U3318 ( .A1(n1750), .A2(\read_value_mux[19][3] ), .A3(n1748), 
        .A4(\read_value_mux[19][2] ), .A5(n2277), .Y(n2280) );
  OA221X1_RVT U3319 ( .A1(search_data[0]), .A2(n1575), .A3(n1752), .A4(
        \read_value_mux[19][0] ), .A5(search), .Y(n2278) );
  OA221X1_RVT U3320 ( .A1(search_data[31]), .A2(n1655), .A3(n1767), .A4(
        \read_value_mux[19][31] ), .A5(n2278), .Y(n2279) );
  NAND4X0_RVT U3321 ( .A1(n2282), .A2(n2281), .A3(n2280), .A4(n2279), .Y(n2283) );
  AO22X1_RVT U3322 ( .A1(search_data[28]), .A2(\read_value_mux[21][28] ), .A3(
        n1758), .A4(n1561), .Y(n2287) );
  OA221X1_RVT U3323 ( .A1(search_data[1]), .A2(n66), .A3(n1755), .A4(
        \read_value_mux[21][1] ), .A5(n2287), .Y(n2294) );
  AO22X1_RVT U3324 ( .A1(search_data[30]), .A2(\read_value_mux[21][30] ), .A3(
        n1764), .A4(n67), .Y(n2288) );
  OA221X1_RVT U3325 ( .A1(search_data[29]), .A2(n1609), .A3(n1761), .A4(
        \read_value_mux[21][29] ), .A5(n2288), .Y(n2293) );
  AOI22X1_RVT U3326 ( .A1(n1543), .A2(\read_value_mux[21][26] ), .A3(n1542), 
        .A4(\read_value_mux[21][27] ), .Y(n2289) );
  OA221X1_RVT U3327 ( .A1(n1542), .A2(\read_value_mux[21][27] ), .A3(n1692), 
        .A4(\read_value_mux[21][26] ), .A5(n2289), .Y(n2292) );
  AOI22X1_RVT U3328 ( .A1(n1541), .A2(\read_value_mux[21][24] ), .A3(n1540), 
        .A4(\read_value_mux[21][25] ), .Y(n2290) );
  OA221X1_RVT U3329 ( .A1(n1540), .A2(\read_value_mux[21][25] ), .A3(n1696), 
        .A4(\read_value_mux[21][24] ), .A5(n2290), .Y(n2291) );
  NAND4X0_RVT U3330 ( .A1(n2294), .A2(n2293), .A3(n2292), .A4(n2291), .Y(n2322) );
  AOI22X1_RVT U3331 ( .A1(n1539), .A2(\read_value_mux[21][22] ), .A3(n1538), 
        .A4(\read_value_mux[21][23] ), .Y(n2295) );
  OA221X1_RVT U3332 ( .A1(n1538), .A2(\read_value_mux[21][23] ), .A3(n1699), 
        .A4(\read_value_mux[21][22] ), .A5(n2295), .Y(n2302) );
  AOI22X1_RVT U3333 ( .A1(n1537), .A2(\read_value_mux[21][20] ), .A3(n1536), 
        .A4(\read_value_mux[21][21] ), .Y(n2296) );
  OA221X1_RVT U3334 ( .A1(n1703), .A2(\read_value_mux[21][21] ), .A3(n1702), 
        .A4(\read_value_mux[21][20] ), .A5(n2296), .Y(n2301) );
  AOI22X1_RVT U3335 ( .A1(n1535), .A2(\read_value_mux[21][18] ), .A3(n1534), 
        .A4(\read_value_mux[21][19] ), .Y(n2297) );
  OA221X1_RVT U3336 ( .A1(n1708), .A2(\read_value_mux[21][19] ), .A3(n1706), 
        .A4(\read_value_mux[21][18] ), .A5(n2297), .Y(n2300) );
  AOI22X1_RVT U3337 ( .A1(n1533), .A2(\read_value_mux[21][16] ), .A3(n1712), 
        .A4(\read_value_mux[21][17] ), .Y(n2298) );
  OA221X1_RVT U3338 ( .A1(n1714), .A2(\read_value_mux[21][17] ), .A3(n1711), 
        .A4(\read_value_mux[21][16] ), .A5(n2298), .Y(n2299) );
  NAND4X0_RVT U3339 ( .A1(n2302), .A2(n2301), .A3(n2300), .A4(n2299), .Y(n2321) );
  AOI22X1_RVT U3340 ( .A1(n1532), .A2(\read_value_mux[21][14] ), .A3(n1719), 
        .A4(\read_value_mux[21][15] ), .Y(n2303) );
  OA221X1_RVT U3341 ( .A1(n1721), .A2(\read_value_mux[21][15] ), .A3(n1717), 
        .A4(\read_value_mux[21][14] ), .A5(n2303), .Y(n2310) );
  AOI22X1_RVT U3342 ( .A1(n1531), .A2(\read_value_mux[21][12] ), .A3(n1530), 
        .A4(\read_value_mux[21][13] ), .Y(n2304) );
  OA221X1_RVT U3343 ( .A1(n1530), .A2(\read_value_mux[21][13] ), .A3(n1725), 
        .A4(\read_value_mux[21][12] ), .A5(n2304), .Y(n2309) );
  AOI22X1_RVT U3344 ( .A1(n1529), .A2(\read_value_mux[21][10] ), .A3(n1528), 
        .A4(\read_value_mux[21][11] ), .Y(n2305) );
  OA221X1_RVT U3345 ( .A1(n1730), .A2(\read_value_mux[21][11] ), .A3(n1728), 
        .A4(\read_value_mux[21][10] ), .A5(n2305), .Y(n2308) );
  AOI22X1_RVT U3346 ( .A1(n1527), .A2(\read_value_mux[21][8] ), .A3(n1734), 
        .A4(\read_value_mux[21][9] ), .Y(n2306) );
  OA221X1_RVT U3347 ( .A1(n1736), .A2(\read_value_mux[21][9] ), .A3(n1733), 
        .A4(\read_value_mux[21][8] ), .A5(n2306), .Y(n2307) );
  NAND4X0_RVT U3348 ( .A1(n2310), .A2(n2309), .A3(n2308), .A4(n2307), .Y(n2320) );
  AOI22X1_RVT U3349 ( .A1(n2940), .A2(\read_value_mux[21][6] ), .A3(n1741), 
        .A4(\read_value_mux[21][7] ), .Y(n2311) );
  OA221X1_RVT U3350 ( .A1(n1740), .A2(\read_value_mux[21][7] ), .A3(n1738), 
        .A4(\read_value_mux[21][6] ), .A5(n2311), .Y(n2318) );
  AOI22X1_RVT U3351 ( .A1(n1526), .A2(\read_value_mux[21][4] ), .A3(n1525), 
        .A4(\read_value_mux[21][5] ), .Y(n2312) );
  OA221X1_RVT U3352 ( .A1(n1745), .A2(\read_value_mux[21][5] ), .A3(n1743), 
        .A4(\read_value_mux[21][4] ), .A5(n2312), .Y(n2317) );
  AOI22X1_RVT U3353 ( .A1(n1524), .A2(\read_value_mux[21][2] ), .A3(n1750), 
        .A4(\read_value_mux[21][3] ), .Y(n2313) );
  OA221X1_RVT U3354 ( .A1(n1750), .A2(\read_value_mux[21][3] ), .A3(n1748), 
        .A4(\read_value_mux[21][2] ), .A5(n2313), .Y(n2316) );
  OA221X1_RVT U3355 ( .A1(search_data[0]), .A2(n1610), .A3(n1752), .A4(
        \read_value_mux[21][0] ), .A5(search), .Y(n2314) );
  OA221X1_RVT U3356 ( .A1(search_data[31]), .A2(n1611), .A3(n1767), .A4(
        \read_value_mux[21][31] ), .A5(n2314), .Y(n2315) );
  NAND4X0_RVT U3357 ( .A1(n2318), .A2(n2317), .A3(n2316), .A4(n2315), .Y(n2319) );
  AO22X1_RVT U3358 ( .A1(search_data[28]), .A2(\read_value_mux[23][28] ), .A3(
        n1758), .A4(n1548), .Y(n2323) );
  OA221X1_RVT U3359 ( .A1(search_data[1]), .A2(n71), .A3(n1755), .A4(
        \read_value_mux[23][1] ), .A5(n2323), .Y(n2330) );
  AO22X1_RVT U3360 ( .A1(search_data[30]), .A2(\read_value_mux[23][30] ), .A3(
        n1764), .A4(n72), .Y(n2324) );
  OA221X1_RVT U3361 ( .A1(search_data[29]), .A2(n1576), .A3(n1761), .A4(
        \read_value_mux[23][29] ), .A5(n2324), .Y(n2329) );
  AOI22X1_RVT U3362 ( .A1(n1543), .A2(\read_value_mux[23][26] ), .A3(n1542), 
        .A4(\read_value_mux[23][27] ), .Y(n2325) );
  OA221X1_RVT U3363 ( .A1(n1542), .A2(\read_value_mux[23][27] ), .A3(n1692), 
        .A4(\read_value_mux[23][26] ), .A5(n2325), .Y(n2328) );
  AOI22X1_RVT U3364 ( .A1(n1541), .A2(\read_value_mux[23][24] ), .A3(n1540), 
        .A4(\read_value_mux[23][25] ), .Y(n2326) );
  OA221X1_RVT U3365 ( .A1(n1540), .A2(\read_value_mux[23][25] ), .A3(n1696), 
        .A4(\read_value_mux[23][24] ), .A5(n2326), .Y(n2327) );
  NAND4X0_RVT U3366 ( .A1(n2330), .A2(n2329), .A3(n2328), .A4(n2327), .Y(n2358) );
  AOI22X1_RVT U3367 ( .A1(n1539), .A2(\read_value_mux[23][22] ), .A3(n1538), 
        .A4(\read_value_mux[23][23] ), .Y(n2331) );
  OA221X1_RVT U3368 ( .A1(n1538), .A2(\read_value_mux[23][23] ), .A3(n1699), 
        .A4(\read_value_mux[23][22] ), .A5(n2331), .Y(n2338) );
  AOI22X1_RVT U3369 ( .A1(n1537), .A2(\read_value_mux[23][20] ), .A3(n1536), 
        .A4(\read_value_mux[23][21] ), .Y(n2332) );
  OA221X1_RVT U3370 ( .A1(n1536), .A2(\read_value_mux[23][21] ), .A3(n1702), 
        .A4(\read_value_mux[23][20] ), .A5(n2332), .Y(n2337) );
  AOI22X1_RVT U3371 ( .A1(n1535), .A2(\read_value_mux[23][18] ), .A3(n1534), 
        .A4(\read_value_mux[23][19] ), .Y(n2333) );
  OA221X1_RVT U3372 ( .A1(n1534), .A2(\read_value_mux[23][19] ), .A3(n1706), 
        .A4(\read_value_mux[23][18] ), .A5(n2333), .Y(n2336) );
  AOI22X1_RVT U3373 ( .A1(n1533), .A2(\read_value_mux[23][16] ), .A3(n1712), 
        .A4(\read_value_mux[23][17] ), .Y(n2334) );
  OA221X1_RVT U3374 ( .A1(n1712), .A2(\read_value_mux[23][17] ), .A3(n1711), 
        .A4(\read_value_mux[23][16] ), .A5(n2334), .Y(n2335) );
  NAND4X0_RVT U3375 ( .A1(n2338), .A2(n2337), .A3(n2336), .A4(n2335), .Y(n2357) );
  AOI22X1_RVT U3376 ( .A1(n1532), .A2(\read_value_mux[23][14] ), .A3(n1719), 
        .A4(\read_value_mux[23][15] ), .Y(n2339) );
  OA221X1_RVT U3377 ( .A1(n1721), .A2(\read_value_mux[23][15] ), .A3(n1717), 
        .A4(\read_value_mux[23][14] ), .A5(n2339), .Y(n2346) );
  AOI22X1_RVT U3378 ( .A1(n1531), .A2(\read_value_mux[23][12] ), .A3(n1530), 
        .A4(\read_value_mux[23][13] ), .Y(n2340) );
  OA221X1_RVT U3379 ( .A1(n1530), .A2(\read_value_mux[23][13] ), .A3(n1725), 
        .A4(\read_value_mux[23][12] ), .A5(n2340), .Y(n2345) );
  AOI22X1_RVT U3380 ( .A1(n1529), .A2(\read_value_mux[23][10] ), .A3(n1528), 
        .A4(\read_value_mux[23][11] ), .Y(n2341) );
  OA221X1_RVT U3381 ( .A1(n1528), .A2(\read_value_mux[23][11] ), .A3(n1728), 
        .A4(\read_value_mux[23][10] ), .A5(n2341), .Y(n2344) );
  AOI22X1_RVT U3382 ( .A1(n1527), .A2(\read_value_mux[23][8] ), .A3(n1734), 
        .A4(\read_value_mux[23][9] ), .Y(n2342) );
  OA221X1_RVT U3383 ( .A1(n1734), .A2(\read_value_mux[23][9] ), .A3(n1733), 
        .A4(\read_value_mux[23][8] ), .A5(n2342), .Y(n2343) );
  NAND4X0_RVT U3384 ( .A1(n2346), .A2(n2345), .A3(n2344), .A4(n2343), .Y(n2356) );
  AOI22X1_RVT U3385 ( .A1(n1738), .A2(\read_value_mux[23][6] ), .A3(n1739), 
        .A4(\read_value_mux[23][7] ), .Y(n2347) );
  OA221X1_RVT U3386 ( .A1(n1740), .A2(\read_value_mux[23][7] ), .A3(n1738), 
        .A4(\read_value_mux[23][6] ), .A5(n2347), .Y(n2354) );
  AOI22X1_RVT U3387 ( .A1(n1526), .A2(\read_value_mux[23][4] ), .A3(n1525), 
        .A4(\read_value_mux[23][5] ), .Y(n2348) );
  OA221X1_RVT U3388 ( .A1(n1745), .A2(\read_value_mux[23][5] ), .A3(n1743), 
        .A4(\read_value_mux[23][4] ), .A5(n2348), .Y(n2353) );
  AOI22X1_RVT U3389 ( .A1(n1524), .A2(\read_value_mux[23][2] ), .A3(n1750), 
        .A4(\read_value_mux[23][3] ), .Y(n2349) );
  OA221X1_RVT U3390 ( .A1(n1750), .A2(\read_value_mux[23][3] ), .A3(n1748), 
        .A4(\read_value_mux[23][2] ), .A5(n2349), .Y(n2352) );
  OA221X1_RVT U3391 ( .A1(search_data[0]), .A2(n1577), .A3(n1752), .A4(
        \read_value_mux[23][0] ), .A5(search), .Y(n2350) );
  OA221X1_RVT U3392 ( .A1(search_data[31]), .A2(n1578), .A3(n1767), .A4(
        \read_value_mux[23][31] ), .A5(n2350), .Y(n2351) );
  NAND4X0_RVT U3393 ( .A1(n2354), .A2(n2353), .A3(n2352), .A4(n2351), .Y(n2355) );
  AO22X1_RVT U3394 ( .A1(search_data[28]), .A2(\read_value_mux[22][28] ), .A3(
        n1758), .A4(n1562), .Y(n2359) );
  OA221X1_RVT U3395 ( .A1(search_data[1]), .A2(n69), .A3(n1755), .A4(
        \read_value_mux[22][1] ), .A5(n2359), .Y(n2366) );
  AO22X1_RVT U3396 ( .A1(search_data[30]), .A2(\read_value_mux[22][30] ), .A3(
        n1764), .A4(n70), .Y(n2360) );
  OA221X1_RVT U3397 ( .A1(search_data[29]), .A2(n1612), .A3(n1761), .A4(
        \read_value_mux[22][29] ), .A5(n2360), .Y(n2365) );
  AOI22X1_RVT U3398 ( .A1(n1691), .A2(\read_value_mux[22][26] ), .A3(n1542), 
        .A4(\read_value_mux[22][27] ), .Y(n2361) );
  OA221X1_RVT U3399 ( .A1(n1542), .A2(\read_value_mux[22][27] ), .A3(n1692), 
        .A4(\read_value_mux[22][26] ), .A5(n2361), .Y(n2364) );
  AOI22X1_RVT U3400 ( .A1(n1695), .A2(\read_value_mux[22][24] ), .A3(n1540), 
        .A4(\read_value_mux[22][25] ), .Y(n2362) );
  OA221X1_RVT U3401 ( .A1(n1540), .A2(\read_value_mux[22][25] ), .A3(n1696), 
        .A4(\read_value_mux[22][24] ), .A5(n2362), .Y(n2363) );
  NAND4X0_RVT U3402 ( .A1(n2366), .A2(n2365), .A3(n2364), .A4(n2363), .Y(n2394) );
  AOI22X1_RVT U3403 ( .A1(n1698), .A2(\read_value_mux[22][22] ), .A3(n1538), 
        .A4(\read_value_mux[22][23] ), .Y(n2367) );
  OA221X1_RVT U3404 ( .A1(n1538), .A2(\read_value_mux[22][23] ), .A3(n1699), 
        .A4(\read_value_mux[22][22] ), .A5(n2367), .Y(n2374) );
  AOI22X1_RVT U3405 ( .A1(n1701), .A2(\read_value_mux[22][20] ), .A3(n1536), 
        .A4(\read_value_mux[22][21] ), .Y(n2368) );
  OA221X1_RVT U3406 ( .A1(n1703), .A2(\read_value_mux[22][21] ), .A3(n1702), 
        .A4(\read_value_mux[22][20] ), .A5(n2368), .Y(n2373) );
  AOI22X1_RVT U3407 ( .A1(n1705), .A2(\read_value_mux[22][18] ), .A3(n1534), 
        .A4(\read_value_mux[22][19] ), .Y(n2369) );
  OA221X1_RVT U3408 ( .A1(n1708), .A2(\read_value_mux[22][19] ), .A3(n1706), 
        .A4(\read_value_mux[22][18] ), .A5(n2369), .Y(n2372) );
  AOI22X1_RVT U3409 ( .A1(n1710), .A2(\read_value_mux[22][16] ), .A3(n1712), 
        .A4(\read_value_mux[22][17] ), .Y(n2370) );
  OA221X1_RVT U3410 ( .A1(n1714), .A2(\read_value_mux[22][17] ), .A3(n1711), 
        .A4(\read_value_mux[22][16] ), .A5(n2370), .Y(n2371) );
  NAND4X0_RVT U3411 ( .A1(n2374), .A2(n2373), .A3(n2372), .A4(n2371), .Y(n2393) );
  AOI22X1_RVT U3412 ( .A1(n1716), .A2(\read_value_mux[22][14] ), .A3(n1719), 
        .A4(\read_value_mux[22][15] ), .Y(n2375) );
  OA221X1_RVT U3413 ( .A1(n1721), .A2(\read_value_mux[22][15] ), .A3(n1717), 
        .A4(\read_value_mux[22][14] ), .A5(n2375), .Y(n2382) );
  AOI22X1_RVT U3414 ( .A1(n1724), .A2(\read_value_mux[22][12] ), .A3(n1530), 
        .A4(\read_value_mux[22][13] ), .Y(n2376) );
  OA221X1_RVT U3415 ( .A1(n1530), .A2(\read_value_mux[22][13] ), .A3(n1725), 
        .A4(\read_value_mux[22][12] ), .A5(n2376), .Y(n2381) );
  AOI22X1_RVT U3416 ( .A1(n1727), .A2(\read_value_mux[22][10] ), .A3(n1528), 
        .A4(\read_value_mux[22][11] ), .Y(n2377) );
  OA221X1_RVT U3417 ( .A1(n1730), .A2(\read_value_mux[22][11] ), .A3(n1728), 
        .A4(\read_value_mux[22][10] ), .A5(n2377), .Y(n2380) );
  AOI22X1_RVT U3418 ( .A1(n1732), .A2(\read_value_mux[22][8] ), .A3(n1734), 
        .A4(\read_value_mux[22][9] ), .Y(n2378) );
  OA221X1_RVT U3419 ( .A1(n1736), .A2(\read_value_mux[22][9] ), .A3(n1733), 
        .A4(\read_value_mux[22][8] ), .A5(n2378), .Y(n2379) );
  NAND4X0_RVT U3420 ( .A1(n2382), .A2(n2381), .A3(n2380), .A4(n2379), .Y(n2392) );
  AOI22X1_RVT U3421 ( .A1(n2940), .A2(\read_value_mux[22][6] ), .A3(n1741), 
        .A4(\read_value_mux[22][7] ), .Y(n2383) );
  OA221X1_RVT U3422 ( .A1(n1740), .A2(\read_value_mux[22][7] ), .A3(n1738), 
        .A4(\read_value_mux[22][6] ), .A5(n2383), .Y(n2390) );
  AOI22X1_RVT U3423 ( .A1(n1742), .A2(\read_value_mux[22][4] ), .A3(n1525), 
        .A4(\read_value_mux[22][5] ), .Y(n2384) );
  OA221X1_RVT U3424 ( .A1(n1745), .A2(\read_value_mux[22][5] ), .A3(n1743), 
        .A4(\read_value_mux[22][4] ), .A5(n2384), .Y(n2389) );
  AOI22X1_RVT U3425 ( .A1(n1524), .A2(\read_value_mux[22][2] ), .A3(n1750), 
        .A4(\read_value_mux[22][3] ), .Y(n2385) );
  OA221X1_RVT U3426 ( .A1(n1750), .A2(\read_value_mux[22][3] ), .A3(n1748), 
        .A4(\read_value_mux[22][2] ), .A5(n2385), .Y(n2388) );
  OA221X1_RVT U3427 ( .A1(search_data[0]), .A2(n1613), .A3(n1752), .A4(
        \read_value_mux[22][0] ), .A5(search), .Y(n2386) );
  OA221X1_RVT U3428 ( .A1(search_data[31]), .A2(n1614), .A3(n1767), .A4(
        \read_value_mux[22][31] ), .A5(n2386), .Y(n2387) );
  NAND4X0_RVT U3429 ( .A1(n2390), .A2(n2389), .A3(n2388), .A4(n2387), .Y(n2391) );
  AO22X1_RVT U3430 ( .A1(search_data[28]), .A2(\read_value_mux[20][28] ), .A3(
        n1758), .A4(n1549), .Y(n2395) );
  OA221X1_RVT U3431 ( .A1(search_data[1]), .A2(n64), .A3(n1755), .A4(
        \read_value_mux[20][1] ), .A5(n2395), .Y(n2402) );
  AO22X1_RVT U3432 ( .A1(search_data[30]), .A2(\read_value_mux[20][30] ), .A3(
        n1764), .A4(n65), .Y(n2396) );
  OA221X1_RVT U3433 ( .A1(search_data[29]), .A2(n1579), .A3(n1761), .A4(
        \read_value_mux[20][29] ), .A5(n2396), .Y(n2401) );
  AOI22X1_RVT U3434 ( .A1(n1691), .A2(\read_value_mux[20][26] ), .A3(n1542), 
        .A4(\read_value_mux[20][27] ), .Y(n2397) );
  OA221X1_RVT U3435 ( .A1(n1542), .A2(\read_value_mux[20][27] ), .A3(n1692), 
        .A4(\read_value_mux[20][26] ), .A5(n2397), .Y(n2400) );
  AOI22X1_RVT U3436 ( .A1(n1695), .A2(\read_value_mux[20][24] ), .A3(n1540), 
        .A4(\read_value_mux[20][25] ), .Y(n2398) );
  OA221X1_RVT U3437 ( .A1(n1540), .A2(\read_value_mux[20][25] ), .A3(n1696), 
        .A4(\read_value_mux[20][24] ), .A5(n2398), .Y(n2399) );
  NAND4X0_RVT U3438 ( .A1(n2402), .A2(n2401), .A3(n2400), .A4(n2399), .Y(n2430) );
  AOI22X1_RVT U3439 ( .A1(n1698), .A2(\read_value_mux[20][22] ), .A3(n1538), 
        .A4(\read_value_mux[20][23] ), .Y(n2403) );
  OA221X1_RVT U3440 ( .A1(n1538), .A2(\read_value_mux[20][23] ), .A3(n1699), 
        .A4(\read_value_mux[20][22] ), .A5(n2403), .Y(n2410) );
  AOI22X1_RVT U3441 ( .A1(n1701), .A2(\read_value_mux[20][20] ), .A3(n1536), 
        .A4(\read_value_mux[20][21] ), .Y(n2404) );
  OA221X1_RVT U3442 ( .A1(n1703), .A2(\read_value_mux[20][21] ), .A3(n1702), 
        .A4(\read_value_mux[20][20] ), .A5(n2404), .Y(n2409) );
  AOI22X1_RVT U3443 ( .A1(n1705), .A2(\read_value_mux[20][18] ), .A3(n1534), 
        .A4(\read_value_mux[20][19] ), .Y(n2405) );
  OA221X1_RVT U3444 ( .A1(n1708), .A2(\read_value_mux[20][19] ), .A3(n1706), 
        .A4(\read_value_mux[20][18] ), .A5(n2405), .Y(n2408) );
  AOI22X1_RVT U3445 ( .A1(n1710), .A2(\read_value_mux[20][16] ), .A3(n1712), 
        .A4(\read_value_mux[20][17] ), .Y(n2406) );
  OA221X1_RVT U3446 ( .A1(n1714), .A2(\read_value_mux[20][17] ), .A3(n1711), 
        .A4(\read_value_mux[20][16] ), .A5(n2406), .Y(n2407) );
  NAND4X0_RVT U3447 ( .A1(n2410), .A2(n2409), .A3(n2408), .A4(n2407), .Y(n2429) );
  AOI22X1_RVT U3448 ( .A1(n1716), .A2(\read_value_mux[20][14] ), .A3(n1719), 
        .A4(\read_value_mux[20][15] ), .Y(n2411) );
  OA221X1_RVT U3449 ( .A1(n1721), .A2(\read_value_mux[20][15] ), .A3(n1717), 
        .A4(\read_value_mux[20][14] ), .A5(n2411), .Y(n2418) );
  AOI22X1_RVT U3450 ( .A1(n1724), .A2(\read_value_mux[20][12] ), .A3(n1530), 
        .A4(\read_value_mux[20][13] ), .Y(n2412) );
  OA221X1_RVT U3451 ( .A1(n1530), .A2(\read_value_mux[20][13] ), .A3(n1725), 
        .A4(\read_value_mux[20][12] ), .A5(n2412), .Y(n2417) );
  AOI22X1_RVT U3452 ( .A1(n1727), .A2(\read_value_mux[20][10] ), .A3(n1528), 
        .A4(\read_value_mux[20][11] ), .Y(n2413) );
  OA221X1_RVT U3453 ( .A1(n1730), .A2(\read_value_mux[20][11] ), .A3(n1728), 
        .A4(\read_value_mux[20][10] ), .A5(n2413), .Y(n2416) );
  AOI22X1_RVT U3454 ( .A1(n1732), .A2(\read_value_mux[20][8] ), .A3(n1734), 
        .A4(\read_value_mux[20][9] ), .Y(n2414) );
  OA221X1_RVT U3455 ( .A1(n1736), .A2(\read_value_mux[20][9] ), .A3(n1733), 
        .A4(\read_value_mux[20][8] ), .A5(n2414), .Y(n2415) );
  NAND4X0_RVT U3456 ( .A1(n2418), .A2(n2417), .A3(n2416), .A4(n2415), .Y(n2428) );
  AOI22X1_RVT U3457 ( .A1(n2940), .A2(\read_value_mux[20][6] ), .A3(n1741), 
        .A4(\read_value_mux[20][7] ), .Y(n2419) );
  OA221X1_RVT U3458 ( .A1(n1740), .A2(\read_value_mux[20][7] ), .A3(n1738), 
        .A4(\read_value_mux[20][6] ), .A5(n2419), .Y(n2426) );
  AOI22X1_RVT U3459 ( .A1(n1742), .A2(\read_value_mux[20][4] ), .A3(n1525), 
        .A4(\read_value_mux[20][5] ), .Y(n2420) );
  OA221X1_RVT U3460 ( .A1(n1745), .A2(\read_value_mux[20][5] ), .A3(n1743), 
        .A4(\read_value_mux[20][4] ), .A5(n2420), .Y(n2425) );
  AOI22X1_RVT U3461 ( .A1(n1524), .A2(\read_value_mux[20][2] ), .A3(n1750), 
        .A4(\read_value_mux[20][3] ), .Y(n2421) );
  OA221X1_RVT U3462 ( .A1(n1750), .A2(\read_value_mux[20][3] ), .A3(n1748), 
        .A4(\read_value_mux[20][2] ), .A5(n2421), .Y(n2424) );
  OA221X1_RVT U3463 ( .A1(search_data[0]), .A2(n1580), .A3(n1752), .A4(
        \read_value_mux[20][0] ), .A5(search), .Y(n2422) );
  OA221X1_RVT U3464 ( .A1(search_data[31]), .A2(n1581), .A3(n1767), .A4(
        \read_value_mux[20][31] ), .A5(n2422), .Y(n2423) );
  NAND4X0_RVT U3465 ( .A1(n2426), .A2(n2425), .A3(n2424), .A4(n2423), .Y(n2427) );
  OA221X1_RVT U3466 ( .A1(n2957), .A2(n2960), .A3(n2957), .A4(n3103), .A5(
        n2431), .Y(n2468) );
  AO22X1_RVT U3467 ( .A1(search_data[28]), .A2(\read_value_mux[15][28] ), .A3(
        n1758), .A4(n1550), .Y(n2432) );
  OA221X1_RVT U3468 ( .A1(search_data[1]), .A2(n50), .A3(n1755), .A4(
        \read_value_mux[15][1] ), .A5(n2432), .Y(n2439) );
  AO22X1_RVT U3469 ( .A1(search_data[30]), .A2(\read_value_mux[15][30] ), .A3(
        n1764), .A4(n51), .Y(n2433) );
  OA221X1_RVT U3470 ( .A1(search_data[29]), .A2(n1582), .A3(n1761), .A4(
        \read_value_mux[15][29] ), .A5(n2433), .Y(n2438) );
  AOI22X1_RVT U3471 ( .A1(n1543), .A2(\read_value_mux[15][26] ), .A3(n1542), 
        .A4(\read_value_mux[15][27] ), .Y(n2434) );
  OA221X1_RVT U3472 ( .A1(n1542), .A2(\read_value_mux[15][27] ), .A3(n1692), 
        .A4(\read_value_mux[15][26] ), .A5(n2434), .Y(n2437) );
  AOI22X1_RVT U3473 ( .A1(n1695), .A2(\read_value_mux[15][24] ), .A3(n1540), 
        .A4(\read_value_mux[15][25] ), .Y(n2435) );
  OA221X1_RVT U3474 ( .A1(n1540), .A2(\read_value_mux[15][25] ), .A3(n1696), 
        .A4(\read_value_mux[15][24] ), .A5(n2435), .Y(n2436) );
  NAND4X0_RVT U3475 ( .A1(n2439), .A2(n2438), .A3(n2437), .A4(n2436), .Y(n2467) );
  AOI22X1_RVT U3476 ( .A1(n1698), .A2(\read_value_mux[15][22] ), .A3(n1538), 
        .A4(\read_value_mux[15][23] ), .Y(n2440) );
  OA221X1_RVT U3477 ( .A1(n1538), .A2(\read_value_mux[15][23] ), .A3(n1699), 
        .A4(\read_value_mux[15][22] ), .A5(n2440), .Y(n2447) );
  AOI22X1_RVT U3478 ( .A1(n1701), .A2(\read_value_mux[15][20] ), .A3(n1536), 
        .A4(\read_value_mux[15][21] ), .Y(n2441) );
  OA221X1_RVT U3479 ( .A1(n1536), .A2(\read_value_mux[15][21] ), .A3(n1702), 
        .A4(\read_value_mux[15][20] ), .A5(n2441), .Y(n2446) );
  AOI22X1_RVT U3480 ( .A1(n1535), .A2(\read_value_mux[15][18] ), .A3(n1534), 
        .A4(\read_value_mux[15][19] ), .Y(n2442) );
  OA221X1_RVT U3481 ( .A1(n1534), .A2(\read_value_mux[15][19] ), .A3(n1706), 
        .A4(\read_value_mux[15][18] ), .A5(n2442), .Y(n2445) );
  AOI22X1_RVT U3482 ( .A1(n1710), .A2(\read_value_mux[15][16] ), .A3(n1712), 
        .A4(\read_value_mux[15][17] ), .Y(n2443) );
  OA221X1_RVT U3483 ( .A1(n1713), .A2(\read_value_mux[15][17] ), .A3(n1711), 
        .A4(\read_value_mux[15][16] ), .A5(n2443), .Y(n2444) );
  NAND4X0_RVT U3484 ( .A1(n2447), .A2(n2446), .A3(n2445), .A4(n2444), .Y(n2466) );
  AOI22X1_RVT U3485 ( .A1(n1716), .A2(\read_value_mux[15][14] ), .A3(n1719), 
        .A4(\read_value_mux[15][15] ), .Y(n2448) );
  OA221X1_RVT U3486 ( .A1(n1720), .A2(\read_value_mux[15][15] ), .A3(n1717), 
        .A4(\read_value_mux[15][14] ), .A5(n2448), .Y(n2455) );
  AOI22X1_RVT U3487 ( .A1(n1724), .A2(\read_value_mux[15][12] ), .A3(n1530), 
        .A4(\read_value_mux[15][13] ), .Y(n2449) );
  OA221X1_RVT U3488 ( .A1(n1530), .A2(\read_value_mux[15][13] ), .A3(n1725), 
        .A4(\read_value_mux[15][12] ), .A5(n2449), .Y(n2454) );
  AOI22X1_RVT U3489 ( .A1(n1529), .A2(\read_value_mux[15][10] ), .A3(n1528), 
        .A4(\read_value_mux[15][11] ), .Y(n2450) );
  OA221X1_RVT U3490 ( .A1(n1528), .A2(\read_value_mux[15][11] ), .A3(n1728), 
        .A4(\read_value_mux[15][10] ), .A5(n2450), .Y(n2453) );
  AOI22X1_RVT U3491 ( .A1(n1732), .A2(\read_value_mux[15][8] ), .A3(n1734), 
        .A4(\read_value_mux[15][9] ), .Y(n2451) );
  OA221X1_RVT U3492 ( .A1(n1735), .A2(\read_value_mux[15][9] ), .A3(n1733), 
        .A4(\read_value_mux[15][8] ), .A5(n2451), .Y(n2452) );
  NAND4X0_RVT U3493 ( .A1(n2455), .A2(n2454), .A3(n2453), .A4(n2452), .Y(n2465) );
  AOI22X1_RVT U3494 ( .A1(n2940), .A2(\read_value_mux[15][6] ), .A3(n1740), 
        .A4(\read_value_mux[15][7] ), .Y(n2456) );
  OA221X1_RVT U3495 ( .A1(n1739), .A2(\read_value_mux[15][7] ), .A3(n1738), 
        .A4(\read_value_mux[15][6] ), .A5(n2456), .Y(n2463) );
  AOI22X1_RVT U3496 ( .A1(n1742), .A2(\read_value_mux[15][4] ), .A3(n1525), 
        .A4(\read_value_mux[15][5] ), .Y(n2457) );
  OA221X1_RVT U3497 ( .A1(n1525), .A2(\read_value_mux[15][5] ), .A3(n1743), 
        .A4(\read_value_mux[15][4] ), .A5(n2457), .Y(n2462) );
  AOI22X1_RVT U3498 ( .A1(n1524), .A2(\read_value_mux[15][2] ), .A3(n1750), 
        .A4(\read_value_mux[15][3] ), .Y(n2458) );
  OA221X1_RVT U3499 ( .A1(n1750), .A2(\read_value_mux[15][3] ), .A3(n1748), 
        .A4(\read_value_mux[15][2] ), .A5(n2458), .Y(n2461) );
  OA221X1_RVT U3500 ( .A1(search_data[0]), .A2(n1583), .A3(n1752), .A4(
        \read_value_mux[15][0] ), .A5(search), .Y(n2459) );
  OA221X1_RVT U3501 ( .A1(search_data[31]), .A2(n1584), .A3(n1767), .A4(
        \read_value_mux[15][31] ), .A5(n2459), .Y(n2460) );
  NAND4X0_RVT U3502 ( .A1(n2463), .A2(n2462), .A3(n2461), .A4(n2460), .Y(n2464) );
  AO221X1_RVT U3503 ( .A1(n2998), .A2(n2979), .A3(n2998), .A4(n2468), .A5(
        n2969), .Y(n2541) );
  AO22X1_RVT U3504 ( .A1(search_data[28]), .A2(\read_value_mux[17][28] ), .A3(
        n1757), .A4(n1642), .Y(n2469) );
  OA221X1_RVT U3505 ( .A1(search_data[1]), .A2(n55), .A3(n1754), .A4(
        \read_value_mux[17][1] ), .A5(n2469), .Y(n2476) );
  AO22X1_RVT U3506 ( .A1(search_data[30]), .A2(\read_value_mux[17][30] ), .A3(
        n1763), .A4(n56), .Y(n2470) );
  OA221X1_RVT U3507 ( .A1(search_data[29]), .A2(n1671), .A3(n1761), .A4(
        \read_value_mux[17][29] ), .A5(n2470), .Y(n2475) );
  AOI22X1_RVT U3508 ( .A1(n1543), .A2(\read_value_mux[17][26] ), .A3(n1542), 
        .A4(\read_value_mux[17][27] ), .Y(n2471) );
  OA221X1_RVT U3509 ( .A1(n1542), .A2(\read_value_mux[17][27] ), .A3(n1692), 
        .A4(\read_value_mux[17][26] ), .A5(n2471), .Y(n2474) );
  AOI22X1_RVT U3510 ( .A1(n1541), .A2(\read_value_mux[17][24] ), .A3(n1540), 
        .A4(\read_value_mux[17][25] ), .Y(n2472) );
  OA221X1_RVT U3511 ( .A1(n1540), .A2(\read_value_mux[17][25] ), .A3(n1696), 
        .A4(\read_value_mux[17][24] ), .A5(n2472), .Y(n2473) );
  NAND4X0_RVT U3512 ( .A1(n2476), .A2(n2475), .A3(n2474), .A4(n2473), .Y(n2504) );
  AOI22X1_RVT U3513 ( .A1(n1698), .A2(\read_value_mux[17][22] ), .A3(n1538), 
        .A4(\read_value_mux[17][23] ), .Y(n2477) );
  OA221X1_RVT U3514 ( .A1(n1538), .A2(\read_value_mux[17][23] ), .A3(n1699), 
        .A4(\read_value_mux[17][22] ), .A5(n2477), .Y(n2484) );
  AOI22X1_RVT U3515 ( .A1(n1702), .A2(\read_value_mux[17][20] ), .A3(n1536), 
        .A4(\read_value_mux[17][21] ), .Y(n2478) );
  OA221X1_RVT U3516 ( .A1(n1536), .A2(\read_value_mux[17][21] ), .A3(n1702), 
        .A4(\read_value_mux[17][20] ), .A5(n2478), .Y(n2483) );
  AOI22X1_RVT U3517 ( .A1(n1706), .A2(\read_value_mux[17][18] ), .A3(n1534), 
        .A4(\read_value_mux[17][19] ), .Y(n2479) );
  OA221X1_RVT U3518 ( .A1(n1534), .A2(\read_value_mux[17][19] ), .A3(n1706), 
        .A4(\read_value_mux[17][18] ), .A5(n2479), .Y(n2482) );
  AOI22X1_RVT U3519 ( .A1(n1711), .A2(\read_value_mux[17][16] ), .A3(n1712), 
        .A4(\read_value_mux[17][17] ), .Y(n2480) );
  OA221X1_RVT U3520 ( .A1(n1712), .A2(\read_value_mux[17][17] ), .A3(n1711), 
        .A4(\read_value_mux[17][16] ), .A5(n2480), .Y(n2481) );
  NAND4X0_RVT U3521 ( .A1(n2484), .A2(n2483), .A3(n2482), .A4(n2481), .Y(n2503) );
  AOI22X1_RVT U3522 ( .A1(n1716), .A2(\read_value_mux[17][14] ), .A3(n1719), 
        .A4(\read_value_mux[17][15] ), .Y(n2485) );
  OA221X1_RVT U3523 ( .A1(n1721), .A2(\read_value_mux[17][15] ), .A3(n1717), 
        .A4(\read_value_mux[17][14] ), .A5(n2485), .Y(n2492) );
  AOI22X1_RVT U3524 ( .A1(n1531), .A2(\read_value_mux[17][12] ), .A3(n1530), 
        .A4(\read_value_mux[17][13] ), .Y(n2486) );
  OA221X1_RVT U3525 ( .A1(n1530), .A2(\read_value_mux[17][13] ), .A3(n1725), 
        .A4(\read_value_mux[17][12] ), .A5(n2486), .Y(n2491) );
  AOI22X1_RVT U3526 ( .A1(n1529), .A2(\read_value_mux[17][10] ), .A3(n1528), 
        .A4(\read_value_mux[17][11] ), .Y(n2487) );
  OA221X1_RVT U3527 ( .A1(n1528), .A2(\read_value_mux[17][11] ), .A3(n1728), 
        .A4(\read_value_mux[17][10] ), .A5(n2487), .Y(n2490) );
  AOI22X1_RVT U3528 ( .A1(n1527), .A2(\read_value_mux[17][8] ), .A3(n1734), 
        .A4(\read_value_mux[17][9] ), .Y(n2488) );
  OA221X1_RVT U3529 ( .A1(n1734), .A2(\read_value_mux[17][9] ), .A3(n1733), 
        .A4(\read_value_mux[17][8] ), .A5(n2488), .Y(n2489) );
  NAND4X0_RVT U3530 ( .A1(n2492), .A2(n2491), .A3(n2490), .A4(n2489), .Y(n2502) );
  AOI22X1_RVT U3531 ( .A1(n2940), .A2(\read_value_mux[17][6] ), .A3(n1741), 
        .A4(\read_value_mux[17][7] ), .Y(n2493) );
  OA221X1_RVT U3532 ( .A1(n1740), .A2(\read_value_mux[17][7] ), .A3(n1738), 
        .A4(\read_value_mux[17][6] ), .A5(n2493), .Y(n2500) );
  AOI22X1_RVT U3533 ( .A1(n1742), .A2(\read_value_mux[17][4] ), .A3(n1525), 
        .A4(\read_value_mux[17][5] ), .Y(n2494) );
  OA221X1_RVT U3534 ( .A1(n1745), .A2(\read_value_mux[17][5] ), .A3(n1743), 
        .A4(\read_value_mux[17][4] ), .A5(n2494), .Y(n2499) );
  AOI22X1_RVT U3535 ( .A1(n1524), .A2(\read_value_mux[17][2] ), .A3(n1750), 
        .A4(\read_value_mux[17][3] ), .Y(n2495) );
  OA221X1_RVT U3536 ( .A1(n1750), .A2(\read_value_mux[17][3] ), .A3(n1748), 
        .A4(\read_value_mux[17][2] ), .A5(n2495), .Y(n2498) );
  OA221X1_RVT U3537 ( .A1(search_data[0]), .A2(n1672), .A3(n1751), .A4(
        \read_value_mux[17][0] ), .A5(search), .Y(n2496) );
  OA221X1_RVT U3538 ( .A1(search_data[31]), .A2(n1673), .A3(n1767), .A4(
        \read_value_mux[17][31] ), .A5(n2496), .Y(n2497) );
  NAND4X0_RVT U3539 ( .A1(n2500), .A2(n2499), .A3(n2498), .A4(n2497), .Y(n2501) );
  AO22X1_RVT U3540 ( .A1(search_data[28]), .A2(\read_value_mux[14][28] ), .A3(
        n1757), .A4(n1563), .Y(n2505) );
  OA221X1_RVT U3541 ( .A1(search_data[1]), .A2(n48), .A3(n1754), .A4(
        \read_value_mux[14][1] ), .A5(n2505), .Y(n2512) );
  AO22X1_RVT U3542 ( .A1(search_data[30]), .A2(\read_value_mux[14][30] ), .A3(
        n1763), .A4(n49), .Y(n2506) );
  OA221X1_RVT U3543 ( .A1(search_data[29]), .A2(n1615), .A3(n1761), .A4(
        \read_value_mux[14][29] ), .A5(n2506), .Y(n2511) );
  AOI22X1_RVT U3544 ( .A1(n1692), .A2(\read_value_mux[14][26] ), .A3(n1542), 
        .A4(\read_value_mux[14][27] ), .Y(n2507) );
  OA221X1_RVT U3545 ( .A1(n1542), .A2(\read_value_mux[14][27] ), .A3(n1692), 
        .A4(\read_value_mux[14][26] ), .A5(n2507), .Y(n2510) );
  AOI22X1_RVT U3546 ( .A1(n1695), .A2(\read_value_mux[14][24] ), .A3(n1540), 
        .A4(\read_value_mux[14][25] ), .Y(n2508) );
  OA221X1_RVT U3547 ( .A1(n1540), .A2(\read_value_mux[14][25] ), .A3(n1696), 
        .A4(\read_value_mux[14][24] ), .A5(n2508), .Y(n2509) );
  NAND4X0_RVT U3548 ( .A1(n2512), .A2(n2511), .A3(n2510), .A4(n2509), .Y(n2540) );
  AOI22X1_RVT U3549 ( .A1(n1539), .A2(\read_value_mux[14][22] ), .A3(n1538), 
        .A4(\read_value_mux[14][23] ), .Y(n2513) );
  OA221X1_RVT U3550 ( .A1(n1538), .A2(\read_value_mux[14][23] ), .A3(n1699), 
        .A4(\read_value_mux[14][22] ), .A5(n2513), .Y(n2520) );
  AOI22X1_RVT U3551 ( .A1(n1537), .A2(\read_value_mux[14][20] ), .A3(n1536), 
        .A4(\read_value_mux[14][21] ), .Y(n2514) );
  OA221X1_RVT U3552 ( .A1(n1536), .A2(\read_value_mux[14][21] ), .A3(n1702), 
        .A4(\read_value_mux[14][20] ), .A5(n2514), .Y(n2519) );
  AOI22X1_RVT U3553 ( .A1(n1535), .A2(\read_value_mux[14][18] ), .A3(n1534), 
        .A4(\read_value_mux[14][19] ), .Y(n2515) );
  OA221X1_RVT U3554 ( .A1(n1534), .A2(\read_value_mux[14][19] ), .A3(n1706), 
        .A4(\read_value_mux[14][18] ), .A5(n2515), .Y(n2518) );
  AOI22X1_RVT U3555 ( .A1(n1710), .A2(\read_value_mux[14][16] ), .A3(n1712), 
        .A4(\read_value_mux[14][17] ), .Y(n2516) );
  OA221X1_RVT U3556 ( .A1(n1713), .A2(\read_value_mux[14][17] ), .A3(n1711), 
        .A4(\read_value_mux[14][16] ), .A5(n2516), .Y(n2517) );
  NAND4X0_RVT U3557 ( .A1(n2520), .A2(n2519), .A3(n2518), .A4(n2517), .Y(n2539) );
  AOI22X1_RVT U3558 ( .A1(n1532), .A2(\read_value_mux[14][14] ), .A3(n1719), 
        .A4(\read_value_mux[14][15] ), .Y(n2521) );
  OA221X1_RVT U3559 ( .A1(n1720), .A2(\read_value_mux[14][15] ), .A3(n1717), 
        .A4(\read_value_mux[14][14] ), .A5(n2521), .Y(n2528) );
  AOI22X1_RVT U3560 ( .A1(n1724), .A2(\read_value_mux[14][12] ), .A3(n1530), 
        .A4(\read_value_mux[14][13] ), .Y(n2522) );
  OA221X1_RVT U3561 ( .A1(n1530), .A2(\read_value_mux[14][13] ), .A3(n1725), 
        .A4(\read_value_mux[14][12] ), .A5(n2522), .Y(n2527) );
  AOI22X1_RVT U3562 ( .A1(n1728), .A2(\read_value_mux[14][10] ), .A3(n1528), 
        .A4(\read_value_mux[14][11] ), .Y(n2523) );
  OA221X1_RVT U3563 ( .A1(n1528), .A2(\read_value_mux[14][11] ), .A3(n1728), 
        .A4(\read_value_mux[14][10] ), .A5(n2523), .Y(n2526) );
  AOI22X1_RVT U3564 ( .A1(n1732), .A2(\read_value_mux[14][8] ), .A3(n1734), 
        .A4(\read_value_mux[14][9] ), .Y(n2524) );
  OA221X1_RVT U3565 ( .A1(n1735), .A2(\read_value_mux[14][9] ), .A3(n1733), 
        .A4(\read_value_mux[14][8] ), .A5(n2524), .Y(n2525) );
  NAND4X0_RVT U3566 ( .A1(n2528), .A2(n2527), .A3(n2526), .A4(n2525), .Y(n2538) );
  AOI22X1_RVT U3567 ( .A1(n2940), .A2(\read_value_mux[14][6] ), .A3(n1741), 
        .A4(\read_value_mux[14][7] ), .Y(n2529) );
  OA221X1_RVT U3568 ( .A1(n1739), .A2(\read_value_mux[14][7] ), .A3(n1738), 
        .A4(\read_value_mux[14][6] ), .A5(n2529), .Y(n2536) );
  AOI22X1_RVT U3569 ( .A1(n1526), .A2(\read_value_mux[14][4] ), .A3(n1525), 
        .A4(\read_value_mux[14][5] ), .Y(n2530) );
  OA221X1_RVT U3570 ( .A1(n1525), .A2(\read_value_mux[14][5] ), .A3(n1743), 
        .A4(\read_value_mux[14][4] ), .A5(n2530), .Y(n2535) );
  AOI22X1_RVT U3571 ( .A1(n1524), .A2(\read_value_mux[14][2] ), .A3(n1750), 
        .A4(\read_value_mux[14][3] ), .Y(n2531) );
  OA221X1_RVT U3572 ( .A1(n1750), .A2(\read_value_mux[14][3] ), .A3(n1748), 
        .A4(\read_value_mux[14][2] ), .A5(n2531), .Y(n2534) );
  OA221X1_RVT U3573 ( .A1(search_data[0]), .A2(n1616), .A3(n1751), .A4(
        \read_value_mux[14][0] ), .A5(search), .Y(n2532) );
  OA221X1_RVT U3574 ( .A1(search_data[31]), .A2(n1617), .A3(n1767), .A4(
        \read_value_mux[14][31] ), .A5(n2532), .Y(n2533) );
  NAND4X0_RVT U3575 ( .A1(n2536), .A2(n2535), .A3(n2534), .A4(n2533), .Y(n2537) );
  OA221X1_RVT U3576 ( .A1(n2541), .A2(n2959), .A3(n2541), .A4(n2985), .A5(
        n2971), .Y(n2578) );
  AO22X1_RVT U3577 ( .A1(search_data[28]), .A2(\read_value_mux[11][28] ), .A3(
        n1757), .A4(n1551), .Y(n2542) );
  OA221X1_RVT U3578 ( .A1(search_data[1]), .A2(n39), .A3(n1754), .A4(
        \read_value_mux[11][1] ), .A5(n2542), .Y(n2549) );
  AO22X1_RVT U3579 ( .A1(search_data[30]), .A2(\read_value_mux[11][30] ), .A3(
        n1763), .A4(n40), .Y(n2543) );
  OA221X1_RVT U3580 ( .A1(search_data[29]), .A2(n1585), .A3(n1760), .A4(
        \read_value_mux[11][29] ), .A5(n2543), .Y(n2548) );
  AOI22X1_RVT U3581 ( .A1(n1691), .A2(\read_value_mux[11][26] ), .A3(n1542), 
        .A4(\read_value_mux[11][27] ), .Y(n2544) );
  OA221X1_RVT U3582 ( .A1(n1542), .A2(\read_value_mux[11][27] ), .A3(n1692), 
        .A4(\read_value_mux[11][26] ), .A5(n2544), .Y(n2547) );
  AOI22X1_RVT U3583 ( .A1(n1541), .A2(\read_value_mux[11][24] ), .A3(n1540), 
        .A4(\read_value_mux[11][25] ), .Y(n2545) );
  OA221X1_RVT U3584 ( .A1(n1540), .A2(\read_value_mux[11][25] ), .A3(n1696), 
        .A4(\read_value_mux[11][24] ), .A5(n2545), .Y(n2546) );
  NAND4X0_RVT U3585 ( .A1(n2549), .A2(n2548), .A3(n2547), .A4(n2546), .Y(n2577) );
  AOI22X1_RVT U3586 ( .A1(n1539), .A2(\read_value_mux[11][22] ), .A3(n1538), 
        .A4(\read_value_mux[11][23] ), .Y(n2550) );
  OA221X1_RVT U3587 ( .A1(n1538), .A2(\read_value_mux[11][23] ), .A3(n1699), 
        .A4(\read_value_mux[11][22] ), .A5(n2550), .Y(n2557) );
  AOI22X1_RVT U3588 ( .A1(n1701), .A2(\read_value_mux[11][20] ), .A3(n1536), 
        .A4(\read_value_mux[11][21] ), .Y(n2551) );
  OA221X1_RVT U3589 ( .A1(n1536), .A2(\read_value_mux[11][21] ), .A3(n1702), 
        .A4(\read_value_mux[11][20] ), .A5(n2551), .Y(n2556) );
  AOI22X1_RVT U3590 ( .A1(n1705), .A2(\read_value_mux[11][18] ), .A3(n1534), 
        .A4(\read_value_mux[11][19] ), .Y(n2552) );
  OA221X1_RVT U3591 ( .A1(n1534), .A2(\read_value_mux[11][19] ), .A3(n1706), 
        .A4(\read_value_mux[11][18] ), .A5(n2552), .Y(n2555) );
  AOI22X1_RVT U3592 ( .A1(n1533), .A2(\read_value_mux[11][16] ), .A3(n1712), 
        .A4(\read_value_mux[11][17] ), .Y(n2553) );
  OA221X1_RVT U3593 ( .A1(n1713), .A2(\read_value_mux[11][17] ), .A3(n1711), 
        .A4(\read_value_mux[11][16] ), .A5(n2553), .Y(n2554) );
  NAND4X0_RVT U3594 ( .A1(n2557), .A2(n2556), .A3(n2555), .A4(n2554), .Y(n2576) );
  AOI22X1_RVT U3595 ( .A1(n1716), .A2(\read_value_mux[11][14] ), .A3(n1719), 
        .A4(\read_value_mux[11][15] ), .Y(n2558) );
  OA221X1_RVT U3596 ( .A1(n1720), .A2(\read_value_mux[11][15] ), .A3(n1717), 
        .A4(\read_value_mux[11][14] ), .A5(n2558), .Y(n2565) );
  AOI22X1_RVT U3597 ( .A1(n1531), .A2(\read_value_mux[11][12] ), .A3(n1530), 
        .A4(\read_value_mux[11][13] ), .Y(n2559) );
  OA221X1_RVT U3598 ( .A1(n1530), .A2(\read_value_mux[11][13] ), .A3(n1725), 
        .A4(\read_value_mux[11][12] ), .A5(n2559), .Y(n2564) );
  AOI22X1_RVT U3599 ( .A1(n1727), .A2(\read_value_mux[11][10] ), .A3(n1528), 
        .A4(\read_value_mux[11][11] ), .Y(n2560) );
  OA221X1_RVT U3600 ( .A1(n1528), .A2(\read_value_mux[11][11] ), .A3(n1728), 
        .A4(\read_value_mux[11][10] ), .A5(n2560), .Y(n2563) );
  AOI22X1_RVT U3601 ( .A1(n1527), .A2(\read_value_mux[11][8] ), .A3(n1734), 
        .A4(\read_value_mux[11][9] ), .Y(n2561) );
  OA221X1_RVT U3602 ( .A1(n1735), .A2(\read_value_mux[11][9] ), .A3(n1733), 
        .A4(\read_value_mux[11][8] ), .A5(n2561), .Y(n2562) );
  NAND4X0_RVT U3603 ( .A1(n2565), .A2(n2564), .A3(n2563), .A4(n2562), .Y(n2575) );
  AOI22X1_RVT U3604 ( .A1(n2940), .A2(\read_value_mux[11][6] ), .A3(n1741), 
        .A4(\read_value_mux[11][7] ), .Y(n2566) );
  OA221X1_RVT U3605 ( .A1(n1739), .A2(\read_value_mux[11][7] ), .A3(n1738), 
        .A4(\read_value_mux[11][6] ), .A5(n2566), .Y(n2573) );
  AOI22X1_RVT U3606 ( .A1(n1526), .A2(\read_value_mux[11][4] ), .A3(n1525), 
        .A4(\read_value_mux[11][5] ), .Y(n2567) );
  OA221X1_RVT U3607 ( .A1(n1525), .A2(\read_value_mux[11][5] ), .A3(n1743), 
        .A4(\read_value_mux[11][4] ), .A5(n2567), .Y(n2572) );
  AOI22X1_RVT U3608 ( .A1(n1524), .A2(\read_value_mux[11][2] ), .A3(n1750), 
        .A4(\read_value_mux[11][3] ), .Y(n2568) );
  OA221X1_RVT U3609 ( .A1(n1750), .A2(\read_value_mux[11][3] ), .A3(n1748), 
        .A4(\read_value_mux[11][2] ), .A5(n2568), .Y(n2571) );
  OA221X1_RVT U3610 ( .A1(search_data[0]), .A2(n1586), .A3(n1751), .A4(
        \read_value_mux[11][0] ), .A5(search), .Y(n2569) );
  OA221X1_RVT U3611 ( .A1(search_data[31]), .A2(n1587), .A3(n1766), .A4(
        \read_value_mux[11][31] ), .A5(n2569), .Y(n2570) );
  NAND4X0_RVT U3612 ( .A1(n2573), .A2(n2572), .A3(n2571), .A4(n2570), .Y(n2574) );
  AO221X1_RVT U3613 ( .A1(n2994), .A2(n2956), .A3(n2994), .A4(n2578), .A5(
        n2973), .Y(n2615) );
  AOI22X1_RVT U3614 ( .A1(n1756), .A2(\read_value_mux[9][1] ), .A3(n1750), 
        .A4(\read_value_mux[9][3] ), .Y(n2579) );
  OA221X1_RVT U3615 ( .A1(n1756), .A2(\read_value_mux[9][1] ), .A3(n1750), 
        .A4(\read_value_mux[9][3] ), .A5(n2579), .Y(n2586) );
  AOI22X1_RVT U3616 ( .A1(n1753), .A2(\read_value_mux[9][0] ), .A3(n1525), 
        .A4(\read_value_mux[9][5] ), .Y(n2580) );
  OA221X1_RVT U3617 ( .A1(n1753), .A2(\read_value_mux[9][0] ), .A3(n1525), 
        .A4(\read_value_mux[9][5] ), .A5(n2580), .Y(n2585) );
  AOI22X1_RVT U3618 ( .A1(n1524), .A2(\read_value_mux[9][2] ), .A3(n1740), 
        .A4(\read_value_mux[9][7] ), .Y(n2581) );
  OA221X1_RVT U3619 ( .A1(n1749), .A2(\read_value_mux[9][2] ), .A3(n1739), 
        .A4(\read_value_mux[9][7] ), .A5(n2581), .Y(n2584) );
  AOI22X1_RVT U3620 ( .A1(n1742), .A2(\read_value_mux[9][4] ), .A3(n1734), 
        .A4(\read_value_mux[9][9] ), .Y(n2582) );
  OA221X1_RVT U3621 ( .A1(n1526), .A2(\read_value_mux[9][4] ), .A3(n1735), 
        .A4(\read_value_mux[9][9] ), .A5(n2582), .Y(n2583) );
  NAND4X0_RVT U3622 ( .A1(n2586), .A2(n2585), .A3(n2584), .A4(n2583), .Y(n2614) );
  AOI22X1_RVT U3623 ( .A1(n2940), .A2(\read_value_mux[9][6] ), .A3(n1528), 
        .A4(\read_value_mux[9][11] ), .Y(n2587) );
  OA221X1_RVT U3624 ( .A1(n2940), .A2(\read_value_mux[9][6] ), .A3(n1528), 
        .A4(\read_value_mux[9][11] ), .A5(n2587), .Y(n2594) );
  AOI22X1_RVT U3625 ( .A1(n1732), .A2(\read_value_mux[9][8] ), .A3(n1530), 
        .A4(\read_value_mux[9][13] ), .Y(n2588) );
  OA221X1_RVT U3626 ( .A1(n1527), .A2(\read_value_mux[9][8] ), .A3(n1530), 
        .A4(\read_value_mux[9][13] ), .A5(n2588), .Y(n2593) );
  AOI22X1_RVT U3627 ( .A1(n1727), .A2(\read_value_mux[9][10] ), .A3(n1719), 
        .A4(\read_value_mux[9][15] ), .Y(n2589) );
  OA221X1_RVT U3628 ( .A1(n1529), .A2(\read_value_mux[9][10] ), .A3(n1720), 
        .A4(\read_value_mux[9][15] ), .A5(n2589), .Y(n2592) );
  AOI22X1_RVT U3629 ( .A1(n1724), .A2(\read_value_mux[9][12] ), .A3(n1712), 
        .A4(\read_value_mux[9][17] ), .Y(n2590) );
  OA221X1_RVT U3630 ( .A1(n1531), .A2(\read_value_mux[9][12] ), .A3(n1713), 
        .A4(\read_value_mux[9][17] ), .A5(n2590), .Y(n2591) );
  NAND4X0_RVT U3631 ( .A1(n2594), .A2(n2593), .A3(n2592), .A4(n2591), .Y(n2613) );
  AOI22X1_RVT U3632 ( .A1(n1716), .A2(\read_value_mux[9][14] ), .A3(n1534), 
        .A4(\read_value_mux[9][19] ), .Y(n2595) );
  OA221X1_RVT U3633 ( .A1(n1532), .A2(\read_value_mux[9][14] ), .A3(n1534), 
        .A4(\read_value_mux[9][19] ), .A5(n2595), .Y(n2602) );
  AOI22X1_RVT U3634 ( .A1(n1710), .A2(\read_value_mux[9][16] ), .A3(n1536), 
        .A4(\read_value_mux[9][21] ), .Y(n2596) );
  OA221X1_RVT U3635 ( .A1(n1533), .A2(\read_value_mux[9][16] ), .A3(n1536), 
        .A4(\read_value_mux[9][21] ), .A5(n2596), .Y(n2601) );
  AOI22X1_RVT U3636 ( .A1(n1705), .A2(\read_value_mux[9][18] ), .A3(n1538), 
        .A4(\read_value_mux[9][23] ), .Y(n2597) );
  OA221X1_RVT U3637 ( .A1(n1535), .A2(\read_value_mux[9][18] ), .A3(n1538), 
        .A4(\read_value_mux[9][23] ), .A5(n2597), .Y(n2600) );
  AOI22X1_RVT U3638 ( .A1(n1701), .A2(\read_value_mux[9][20] ), .A3(n1540), 
        .A4(\read_value_mux[9][25] ), .Y(n2598) );
  OA221X1_RVT U3639 ( .A1(n1537), .A2(\read_value_mux[9][20] ), .A3(n1540), 
        .A4(\read_value_mux[9][25] ), .A5(n2598), .Y(n2599) );
  NAND4X0_RVT U3640 ( .A1(n2602), .A2(n2601), .A3(n2600), .A4(n2599), .Y(n2612) );
  AOI22X1_RVT U3641 ( .A1(n1698), .A2(\read_value_mux[9][22] ), .A3(n1542), 
        .A4(\read_value_mux[9][27] ), .Y(n2603) );
  OA221X1_RVT U3642 ( .A1(n1539), .A2(\read_value_mux[9][22] ), .A3(n1542), 
        .A4(\read_value_mux[9][27] ), .A5(n2603), .Y(n2610) );
  AOI22X1_RVT U3643 ( .A1(n1695), .A2(\read_value_mux[9][24] ), .A3(n1760), 
        .A4(\read_value_mux[9][29] ), .Y(n2604) );
  OA221X1_RVT U3644 ( .A1(n1541), .A2(\read_value_mux[9][24] ), .A3(n1760), 
        .A4(\read_value_mux[9][29] ), .A5(n2604), .Y(n2609) );
  AOI22X1_RVT U3645 ( .A1(n1691), .A2(\read_value_mux[9][26] ), .A3(n1766), 
        .A4(\read_value_mux[9][31] ), .Y(n2605) );
  OA221X1_RVT U3646 ( .A1(n1543), .A2(\read_value_mux[9][26] ), .A3(n1766), 
        .A4(\read_value_mux[9][31] ), .A5(n2605), .Y(n2608) );
  OA221X1_RVT U3647 ( .A1(search_data[28]), .A2(n1618), .A3(n1759), .A4(
        \read_value_mux[9][28] ), .A5(search), .Y(n2606) );
  OA221X1_RVT U3648 ( .A1(search_data[30]), .A2(n34), .A3(n1765), .A4(
        \read_value_mux[9][30] ), .A5(n2606), .Y(n2607) );
  NAND4X0_RVT U3649 ( .A1(n2610), .A2(n2609), .A3(n2608), .A4(n2607), .Y(n2611) );
  AO21X1_RVT U3650 ( .A1(n2975), .A2(n2615), .A3(n2977), .Y(n2955) );
  AO22X1_RVT U3651 ( .A1(search_data[28]), .A2(\read_value_mux[24][28] ), .A3(
        n1757), .A4(n1552), .Y(n2616) );
  OA221X1_RVT U3652 ( .A1(search_data[1]), .A2(n74), .A3(n1754), .A4(
        \read_value_mux[24][1] ), .A5(n2616), .Y(n2623) );
  AO22X1_RVT U3653 ( .A1(search_data[30]), .A2(\read_value_mux[24][30] ), .A3(
        n1763), .A4(n75), .Y(n2617) );
  OA221X1_RVT U3654 ( .A1(search_data[29]), .A2(n1588), .A3(n1760), .A4(
        \read_value_mux[24][29] ), .A5(n2617), .Y(n2622) );
  AOI22X1_RVT U3655 ( .A1(n1543), .A2(\read_value_mux[24][26] ), .A3(n1542), 
        .A4(\read_value_mux[24][27] ), .Y(n2618) );
  OA221X1_RVT U3656 ( .A1(n1542), .A2(\read_value_mux[24][27] ), .A3(n1692), 
        .A4(\read_value_mux[24][26] ), .A5(n2618), .Y(n2621) );
  AOI22X1_RVT U3657 ( .A1(n1541), .A2(\read_value_mux[24][24] ), .A3(n1540), 
        .A4(\read_value_mux[24][25] ), .Y(n2619) );
  OA221X1_RVT U3658 ( .A1(n1540), .A2(\read_value_mux[24][25] ), .A3(n1696), 
        .A4(\read_value_mux[24][24] ), .A5(n2619), .Y(n2620) );
  NAND4X0_RVT U3659 ( .A1(n2623), .A2(n2622), .A3(n2621), .A4(n2620), .Y(n2651) );
  AOI22X1_RVT U3660 ( .A1(n1698), .A2(\read_value_mux[24][22] ), .A3(n1538), 
        .A4(\read_value_mux[24][23] ), .Y(n2624) );
  OA221X1_RVT U3661 ( .A1(n1538), .A2(\read_value_mux[24][23] ), .A3(n1699), 
        .A4(\read_value_mux[24][22] ), .A5(n2624), .Y(n2631) );
  AOI22X1_RVT U3662 ( .A1(n1537), .A2(\read_value_mux[24][20] ), .A3(n1536), 
        .A4(\read_value_mux[24][21] ), .Y(n2625) );
  OA221X1_RVT U3663 ( .A1(n1703), .A2(\read_value_mux[24][21] ), .A3(n1702), 
        .A4(\read_value_mux[24][20] ), .A5(n2625), .Y(n2630) );
  AOI22X1_RVT U3664 ( .A1(n1535), .A2(\read_value_mux[24][18] ), .A3(n1534), 
        .A4(\read_value_mux[24][19] ), .Y(n2626) );
  OA221X1_RVT U3665 ( .A1(n1708), .A2(\read_value_mux[24][19] ), .A3(n1706), 
        .A4(\read_value_mux[24][18] ), .A5(n2626), .Y(n2629) );
  AOI22X1_RVT U3666 ( .A1(n1533), .A2(\read_value_mux[24][16] ), .A3(n1713), 
        .A4(\read_value_mux[24][17] ), .Y(n2627) );
  OA221X1_RVT U3667 ( .A1(n1714), .A2(\read_value_mux[24][17] ), .A3(n1711), 
        .A4(\read_value_mux[24][16] ), .A5(n2627), .Y(n2628) );
  NAND4X0_RVT U3668 ( .A1(n2631), .A2(n2630), .A3(n2629), .A4(n2628), .Y(n2650) );
  AOI22X1_RVT U3669 ( .A1(n1532), .A2(\read_value_mux[24][14] ), .A3(n1720), 
        .A4(\read_value_mux[24][15] ), .Y(n2632) );
  OA221X1_RVT U3670 ( .A1(n1721), .A2(\read_value_mux[24][15] ), .A3(n1717), 
        .A4(\read_value_mux[24][14] ), .A5(n2632), .Y(n2639) );
  AOI22X1_RVT U3671 ( .A1(n1531), .A2(\read_value_mux[24][12] ), .A3(n1530), 
        .A4(\read_value_mux[24][13] ), .Y(n2633) );
  OA221X1_RVT U3672 ( .A1(n1530), .A2(\read_value_mux[24][13] ), .A3(n1725), 
        .A4(\read_value_mux[24][12] ), .A5(n2633), .Y(n2638) );
  AOI22X1_RVT U3673 ( .A1(n1529), .A2(\read_value_mux[24][10] ), .A3(n1528), 
        .A4(\read_value_mux[24][11] ), .Y(n2634) );
  OA221X1_RVT U3674 ( .A1(n1730), .A2(\read_value_mux[24][11] ), .A3(n1728), 
        .A4(\read_value_mux[24][10] ), .A5(n2634), .Y(n2637) );
  AOI22X1_RVT U3675 ( .A1(n1527), .A2(\read_value_mux[24][8] ), .A3(n1735), 
        .A4(\read_value_mux[24][9] ), .Y(n2635) );
  OA221X1_RVT U3676 ( .A1(n1736), .A2(\read_value_mux[24][9] ), .A3(n1733), 
        .A4(\read_value_mux[24][8] ), .A5(n2635), .Y(n2636) );
  NAND4X0_RVT U3677 ( .A1(n2639), .A2(n2638), .A3(n2637), .A4(n2636), .Y(n2649) );
  AOI22X1_RVT U3678 ( .A1(n2940), .A2(\read_value_mux[24][6] ), .A3(n1739), 
        .A4(\read_value_mux[24][7] ), .Y(n2640) );
  OA221X1_RVT U3679 ( .A1(n1740), .A2(\read_value_mux[24][7] ), .A3(n1738), 
        .A4(\read_value_mux[24][6] ), .A5(n2640), .Y(n2647) );
  AOI22X1_RVT U3680 ( .A1(n1742), .A2(\read_value_mux[24][4] ), .A3(n1525), 
        .A4(\read_value_mux[24][5] ), .Y(n2641) );
  OA221X1_RVT U3681 ( .A1(n1745), .A2(\read_value_mux[24][5] ), .A3(n1743), 
        .A4(\read_value_mux[24][4] ), .A5(n2641), .Y(n2646) );
  AOI22X1_RVT U3682 ( .A1(n1524), .A2(\read_value_mux[24][2] ), .A3(n1750), 
        .A4(\read_value_mux[24][3] ), .Y(n2642) );
  OA221X1_RVT U3683 ( .A1(n1750), .A2(\read_value_mux[24][3] ), .A3(n1748), 
        .A4(\read_value_mux[24][2] ), .A5(n2642), .Y(n2645) );
  OA221X1_RVT U3684 ( .A1(search_data[0]), .A2(n1589), .A3(n1751), .A4(
        \read_value_mux[24][0] ), .A5(search), .Y(n2643) );
  OA221X1_RVT U3685 ( .A1(search_data[31]), .A2(n1590), .A3(n1766), .A4(
        \read_value_mux[24][31] ), .A5(n2643), .Y(n2644) );
  NAND4X0_RVT U3686 ( .A1(n2647), .A2(n2646), .A3(n2645), .A4(n2644), .Y(n2648) );
  NAND4X0_RVT U3687 ( .A1(n2975), .A2(n2994), .A3(n2971), .A4(n2962), .Y(n2652) );
  AO22X1_RVT U3688 ( .A1(search_data[28]), .A2(\read_value_mux[26][28] ), .A3(
        n1757), .A4(n1564), .Y(n2655) );
  OA221X1_RVT U3689 ( .A1(search_data[1]), .A2(n79), .A3(n1754), .A4(
        \read_value_mux[26][1] ), .A5(n2655), .Y(n2662) );
  AO22X1_RVT U3690 ( .A1(search_data[30]), .A2(\read_value_mux[26][30] ), .A3(
        n1763), .A4(n80), .Y(n2656) );
  OA221X1_RVT U3691 ( .A1(search_data[29]), .A2(n1619), .A3(n1760), .A4(
        \read_value_mux[26][29] ), .A5(n2656), .Y(n2661) );
  AOI22X1_RVT U3692 ( .A1(n1543), .A2(\read_value_mux[26][26] ), .A3(n1542), 
        .A4(\read_value_mux[26][27] ), .Y(n2657) );
  OA221X1_RVT U3693 ( .A1(n1542), .A2(\read_value_mux[26][27] ), .A3(n1692), 
        .A4(\read_value_mux[26][26] ), .A5(n2657), .Y(n2660) );
  AOI22X1_RVT U3694 ( .A1(n1695), .A2(\read_value_mux[26][24] ), .A3(n1540), 
        .A4(\read_value_mux[26][25] ), .Y(n2658) );
  OA221X1_RVT U3695 ( .A1(n1540), .A2(\read_value_mux[26][25] ), .A3(n1696), 
        .A4(\read_value_mux[26][24] ), .A5(n2658), .Y(n2659) );
  NAND4X0_RVT U3696 ( .A1(n2662), .A2(n2661), .A3(n2660), .A4(n2659), .Y(n2690) );
  AOI22X1_RVT U3697 ( .A1(n1539), .A2(\read_value_mux[26][22] ), .A3(n1538), 
        .A4(\read_value_mux[26][23] ), .Y(n2663) );
  OA221X1_RVT U3698 ( .A1(n1538), .A2(\read_value_mux[26][23] ), .A3(n1699), 
        .A4(\read_value_mux[26][22] ), .A5(n2663), .Y(n2670) );
  AOI22X1_RVT U3699 ( .A1(n1701), .A2(\read_value_mux[26][20] ), .A3(n1536), 
        .A4(\read_value_mux[26][21] ), .Y(n2664) );
  OA221X1_RVT U3700 ( .A1(n1703), .A2(\read_value_mux[26][21] ), .A3(n1702), 
        .A4(\read_value_mux[26][20] ), .A5(n2664), .Y(n2669) );
  AOI22X1_RVT U3701 ( .A1(n1535), .A2(\read_value_mux[26][18] ), .A3(n1534), 
        .A4(\read_value_mux[26][19] ), .Y(n2665) );
  OA221X1_RVT U3702 ( .A1(n1708), .A2(\read_value_mux[26][19] ), .A3(n1706), 
        .A4(\read_value_mux[26][18] ), .A5(n2665), .Y(n2668) );
  AOI22X1_RVT U3703 ( .A1(n1710), .A2(\read_value_mux[26][16] ), .A3(n1712), 
        .A4(\read_value_mux[26][17] ), .Y(n2666) );
  OA221X1_RVT U3704 ( .A1(n1714), .A2(\read_value_mux[26][17] ), .A3(n1711), 
        .A4(\read_value_mux[26][16] ), .A5(n2666), .Y(n2667) );
  NAND4X0_RVT U3705 ( .A1(n2670), .A2(n2669), .A3(n2668), .A4(n2667), .Y(n2689) );
  AOI22X1_RVT U3706 ( .A1(n1532), .A2(\read_value_mux[26][14] ), .A3(n1719), 
        .A4(\read_value_mux[26][15] ), .Y(n2671) );
  OA221X1_RVT U3707 ( .A1(n1721), .A2(\read_value_mux[26][15] ), .A3(n1717), 
        .A4(\read_value_mux[26][14] ), .A5(n2671), .Y(n2678) );
  AOI22X1_RVT U3708 ( .A1(n1724), .A2(\read_value_mux[26][12] ), .A3(n1530), 
        .A4(\read_value_mux[26][13] ), .Y(n2672) );
  OA221X1_RVT U3709 ( .A1(n1530), .A2(\read_value_mux[26][13] ), .A3(n1725), 
        .A4(\read_value_mux[26][12] ), .A5(n2672), .Y(n2677) );
  AOI22X1_RVT U3710 ( .A1(n1529), .A2(\read_value_mux[26][10] ), .A3(n1528), 
        .A4(\read_value_mux[26][11] ), .Y(n2673) );
  OA221X1_RVT U3711 ( .A1(n1730), .A2(\read_value_mux[26][11] ), .A3(n1728), 
        .A4(\read_value_mux[26][10] ), .A5(n2673), .Y(n2676) );
  AOI22X1_RVT U3712 ( .A1(n1732), .A2(\read_value_mux[26][8] ), .A3(n1734), 
        .A4(\read_value_mux[26][9] ), .Y(n2674) );
  OA221X1_RVT U3713 ( .A1(n1736), .A2(\read_value_mux[26][9] ), .A3(n1733), 
        .A4(\read_value_mux[26][8] ), .A5(n2674), .Y(n2675) );
  NAND4X0_RVT U3714 ( .A1(n2678), .A2(n2677), .A3(n2676), .A4(n2675), .Y(n2688) );
  AOI22X1_RVT U3715 ( .A1(n2940), .A2(\read_value_mux[26][6] ), .A3(n1741), 
        .A4(\read_value_mux[26][7] ), .Y(n2679) );
  OA221X1_RVT U3716 ( .A1(n1740), .A2(\read_value_mux[26][7] ), .A3(n1738), 
        .A4(\read_value_mux[26][6] ), .A5(n2679), .Y(n2686) );
  AOI22X1_RVT U3717 ( .A1(n1526), .A2(\read_value_mux[26][4] ), .A3(n1525), 
        .A4(\read_value_mux[26][5] ), .Y(n2680) );
  OA221X1_RVT U3718 ( .A1(n1745), .A2(\read_value_mux[26][5] ), .A3(n1743), 
        .A4(\read_value_mux[26][4] ), .A5(n2680), .Y(n2685) );
  AOI22X1_RVT U3719 ( .A1(n1524), .A2(\read_value_mux[26][2] ), .A3(n1750), 
        .A4(\read_value_mux[26][3] ), .Y(n2681) );
  OA221X1_RVT U3720 ( .A1(n1750), .A2(\read_value_mux[26][3] ), .A3(n1748), 
        .A4(\read_value_mux[26][2] ), .A5(n2681), .Y(n2684) );
  OA221X1_RVT U3721 ( .A1(search_data[0]), .A2(n1620), .A3(n1751), .A4(
        \read_value_mux[26][0] ), .A5(search), .Y(n2682) );
  OA221X1_RVT U3722 ( .A1(search_data[31]), .A2(n1621), .A3(n1766), .A4(
        \read_value_mux[26][31] ), .A5(n2682), .Y(n2683) );
  NAND4X0_RVT U3723 ( .A1(n2686), .A2(n2685), .A3(n2684), .A4(n2683), .Y(n2687) );
  AO22X1_RVT U3724 ( .A1(search_data[28]), .A2(\read_value_mux[27][28] ), .A3(
        n1757), .A4(n1553), .Y(n2691) );
  OA221X1_RVT U3725 ( .A1(search_data[1]), .A2(n81), .A3(n1754), .A4(
        \read_value_mux[27][1] ), .A5(n2691), .Y(n2698) );
  AO22X1_RVT U3726 ( .A1(search_data[30]), .A2(\read_value_mux[27][30] ), .A3(
        n1763), .A4(n82), .Y(n2692) );
  OA221X1_RVT U3727 ( .A1(search_data[29]), .A2(n1591), .A3(n1760), .A4(
        \read_value_mux[27][29] ), .A5(n2692), .Y(n2697) );
  AOI22X1_RVT U3728 ( .A1(n1691), .A2(\read_value_mux[27][26] ), .A3(n1542), 
        .A4(\read_value_mux[27][27] ), .Y(n2693) );
  OA221X1_RVT U3729 ( .A1(n1542), .A2(\read_value_mux[27][27] ), .A3(n1692), 
        .A4(\read_value_mux[27][26] ), .A5(n2693), .Y(n2696) );
  AOI22X1_RVT U3730 ( .A1(n1695), .A2(\read_value_mux[27][24] ), .A3(n1540), 
        .A4(\read_value_mux[27][25] ), .Y(n2694) );
  OA221X1_RVT U3731 ( .A1(n1540), .A2(\read_value_mux[27][25] ), .A3(n1696), 
        .A4(\read_value_mux[27][24] ), .A5(n2694), .Y(n2695) );
  NAND4X0_RVT U3732 ( .A1(n2698), .A2(n2697), .A3(n2696), .A4(n2695), .Y(n2726) );
  AOI22X1_RVT U3733 ( .A1(n1698), .A2(\read_value_mux[27][22] ), .A3(n1538), 
        .A4(\read_value_mux[27][23] ), .Y(n2699) );
  OA221X1_RVT U3734 ( .A1(n1538), .A2(\read_value_mux[27][23] ), .A3(n1699), 
        .A4(\read_value_mux[27][22] ), .A5(n2699), .Y(n2706) );
  AOI22X1_RVT U3735 ( .A1(n1701), .A2(\read_value_mux[27][20] ), .A3(n1536), 
        .A4(\read_value_mux[27][21] ), .Y(n2700) );
  OA221X1_RVT U3736 ( .A1(n1703), .A2(\read_value_mux[27][21] ), .A3(n1702), 
        .A4(\read_value_mux[27][20] ), .A5(n2700), .Y(n2705) );
  AOI22X1_RVT U3737 ( .A1(n1705), .A2(\read_value_mux[27][18] ), .A3(n1534), 
        .A4(\read_value_mux[27][19] ), .Y(n2701) );
  OA221X1_RVT U3738 ( .A1(n1708), .A2(\read_value_mux[27][19] ), .A3(n1706), 
        .A4(\read_value_mux[27][18] ), .A5(n2701), .Y(n2704) );
  AOI22X1_RVT U3739 ( .A1(n1710), .A2(\read_value_mux[27][16] ), .A3(n1713), 
        .A4(\read_value_mux[27][17] ), .Y(n2702) );
  OA221X1_RVT U3740 ( .A1(n1714), .A2(\read_value_mux[27][17] ), .A3(n1711), 
        .A4(\read_value_mux[27][16] ), .A5(n2702), .Y(n2703) );
  NAND4X0_RVT U3741 ( .A1(n2706), .A2(n2705), .A3(n2704), .A4(n2703), .Y(n2725) );
  AOI22X1_RVT U3742 ( .A1(n1716), .A2(\read_value_mux[27][14] ), .A3(n1720), 
        .A4(\read_value_mux[27][15] ), .Y(n2707) );
  OA221X1_RVT U3743 ( .A1(n1721), .A2(\read_value_mux[27][15] ), .A3(n1717), 
        .A4(\read_value_mux[27][14] ), .A5(n2707), .Y(n2714) );
  AOI22X1_RVT U3744 ( .A1(n1724), .A2(\read_value_mux[27][12] ), .A3(n1530), 
        .A4(\read_value_mux[27][13] ), .Y(n2708) );
  OA221X1_RVT U3745 ( .A1(n1530), .A2(\read_value_mux[27][13] ), .A3(n1725), 
        .A4(\read_value_mux[27][12] ), .A5(n2708), .Y(n2713) );
  AOI22X1_RVT U3746 ( .A1(n1727), .A2(\read_value_mux[27][10] ), .A3(n1528), 
        .A4(\read_value_mux[27][11] ), .Y(n2709) );
  OA221X1_RVT U3747 ( .A1(n1730), .A2(\read_value_mux[27][11] ), .A3(n1728), 
        .A4(\read_value_mux[27][10] ), .A5(n2709), .Y(n2712) );
  AOI22X1_RVT U3748 ( .A1(n1732), .A2(\read_value_mux[27][8] ), .A3(n1735), 
        .A4(\read_value_mux[27][9] ), .Y(n2710) );
  OA221X1_RVT U3749 ( .A1(n1736), .A2(\read_value_mux[27][9] ), .A3(n1733), 
        .A4(\read_value_mux[27][8] ), .A5(n2710), .Y(n2711) );
  NAND4X0_RVT U3750 ( .A1(n2714), .A2(n2713), .A3(n2712), .A4(n2711), .Y(n2724) );
  AOI22X1_RVT U3751 ( .A1(n2940), .A2(\read_value_mux[27][6] ), .A3(n1739), 
        .A4(\read_value_mux[27][7] ), .Y(n2715) );
  OA221X1_RVT U3752 ( .A1(n1740), .A2(\read_value_mux[27][7] ), .A3(n1738), 
        .A4(\read_value_mux[27][6] ), .A5(n2715), .Y(n2722) );
  AOI22X1_RVT U3753 ( .A1(n1742), .A2(\read_value_mux[27][4] ), .A3(n1525), 
        .A4(\read_value_mux[27][5] ), .Y(n2716) );
  OA221X1_RVT U3754 ( .A1(n1745), .A2(\read_value_mux[27][5] ), .A3(n1743), 
        .A4(\read_value_mux[27][4] ), .A5(n2716), .Y(n2721) );
  AOI22X1_RVT U3755 ( .A1(n1524), .A2(\read_value_mux[27][2] ), .A3(n1750), 
        .A4(\read_value_mux[27][3] ), .Y(n2717) );
  OA221X1_RVT U3756 ( .A1(n1750), .A2(\read_value_mux[27][3] ), .A3(n1748), 
        .A4(\read_value_mux[27][2] ), .A5(n2717), .Y(n2720) );
  OA221X1_RVT U3757 ( .A1(search_data[0]), .A2(n1592), .A3(n1751), .A4(
        \read_value_mux[27][0] ), .A5(search), .Y(n2718) );
  OA221X1_RVT U3758 ( .A1(search_data[31]), .A2(n1593), .A3(n1766), .A4(
        \read_value_mux[27][31] ), .A5(n2718), .Y(n2719) );
  NAND4X0_RVT U3759 ( .A1(n2722), .A2(n2721), .A3(n2720), .A4(n2719), .Y(n2723) );
  AO22X1_RVT U3760 ( .A1(search_data[28]), .A2(\read_value_mux[29][28] ), .A3(
        n1757), .A4(n1565), .Y(n2727) );
  OA221X1_RVT U3761 ( .A1(search_data[1]), .A2(n85), .A3(n1754), .A4(
        \read_value_mux[29][1] ), .A5(n2727), .Y(n2734) );
  AO22X1_RVT U3762 ( .A1(search_data[30]), .A2(\read_value_mux[29][30] ), .A3(
        n1763), .A4(n86), .Y(n2728) );
  OA221X1_RVT U3763 ( .A1(search_data[29]), .A2(n1622), .A3(n1760), .A4(
        \read_value_mux[29][29] ), .A5(n2728), .Y(n2733) );
  AOI22X1_RVT U3764 ( .A1(n1691), .A2(\read_value_mux[29][26] ), .A3(n1542), 
        .A4(\read_value_mux[29][27] ), .Y(n2729) );
  OA221X1_RVT U3765 ( .A1(n1542), .A2(\read_value_mux[29][27] ), .A3(n1691), 
        .A4(\read_value_mux[29][26] ), .A5(n2729), .Y(n2732) );
  AOI22X1_RVT U3766 ( .A1(n1541), .A2(\read_value_mux[29][24] ), .A3(n1540), 
        .A4(\read_value_mux[29][25] ), .Y(n2730) );
  OA221X1_RVT U3767 ( .A1(n1540), .A2(\read_value_mux[29][25] ), .A3(n1695), 
        .A4(\read_value_mux[29][24] ), .A5(n2730), .Y(n2731) );
  NAND4X0_RVT U3768 ( .A1(n2734), .A2(n2733), .A3(n2732), .A4(n2731), .Y(n2762) );
  AOI22X1_RVT U3769 ( .A1(n1698), .A2(\read_value_mux[29][22] ), .A3(n1538), 
        .A4(\read_value_mux[29][23] ), .Y(n2735) );
  OA221X1_RVT U3770 ( .A1(n1538), .A2(\read_value_mux[29][23] ), .A3(n1698), 
        .A4(\read_value_mux[29][22] ), .A5(n2735), .Y(n2742) );
  AOI22X1_RVT U3771 ( .A1(n1537), .A2(\read_value_mux[29][20] ), .A3(n1536), 
        .A4(\read_value_mux[29][21] ), .Y(n2736) );
  OA221X1_RVT U3772 ( .A1(n1703), .A2(\read_value_mux[29][21] ), .A3(n1701), 
        .A4(\read_value_mux[29][20] ), .A5(n2736), .Y(n2741) );
  AOI22X1_RVT U3773 ( .A1(n1705), .A2(\read_value_mux[29][18] ), .A3(n1534), 
        .A4(\read_value_mux[29][19] ), .Y(n2737) );
  OA221X1_RVT U3774 ( .A1(n1708), .A2(\read_value_mux[29][19] ), .A3(n1705), 
        .A4(\read_value_mux[29][18] ), .A5(n2737), .Y(n2740) );
  AOI22X1_RVT U3775 ( .A1(n1533), .A2(\read_value_mux[29][16] ), .A3(n1713), 
        .A4(\read_value_mux[29][17] ), .Y(n2738) );
  OA221X1_RVT U3776 ( .A1(n1714), .A2(\read_value_mux[29][17] ), .A3(n1710), 
        .A4(\read_value_mux[29][16] ), .A5(n2738), .Y(n2739) );
  NAND4X0_RVT U3777 ( .A1(n2742), .A2(n2741), .A3(n2740), .A4(n2739), .Y(n2761) );
  AOI22X1_RVT U3778 ( .A1(n1716), .A2(\read_value_mux[29][14] ), .A3(n1720), 
        .A4(\read_value_mux[29][15] ), .Y(n2743) );
  OA221X1_RVT U3779 ( .A1(n1721), .A2(\read_value_mux[29][15] ), .A3(n1716), 
        .A4(\read_value_mux[29][14] ), .A5(n2743), .Y(n2750) );
  AOI22X1_RVT U3780 ( .A1(n1531), .A2(\read_value_mux[29][12] ), .A3(n1530), 
        .A4(\read_value_mux[29][13] ), .Y(n2744) );
  OA221X1_RVT U3781 ( .A1(n1530), .A2(\read_value_mux[29][13] ), .A3(n1724), 
        .A4(\read_value_mux[29][12] ), .A5(n2744), .Y(n2749) );
  AOI22X1_RVT U3782 ( .A1(n1727), .A2(\read_value_mux[29][10] ), .A3(n1528), 
        .A4(\read_value_mux[29][11] ), .Y(n2745) );
  OA221X1_RVT U3783 ( .A1(n1730), .A2(\read_value_mux[29][11] ), .A3(n1727), 
        .A4(\read_value_mux[29][10] ), .A5(n2745), .Y(n2748) );
  AOI22X1_RVT U3784 ( .A1(n1527), .A2(\read_value_mux[29][8] ), .A3(n1735), 
        .A4(\read_value_mux[29][9] ), .Y(n2746) );
  OA221X1_RVT U3785 ( .A1(n1736), .A2(\read_value_mux[29][9] ), .A3(n1732), 
        .A4(\read_value_mux[29][8] ), .A5(n2746), .Y(n2747) );
  NAND4X0_RVT U3786 ( .A1(n2750), .A2(n2749), .A3(n2748), .A4(n2747), .Y(n2760) );
  AOI22X1_RVT U3787 ( .A1(n2940), .A2(\read_value_mux[29][6] ), .A3(n1739), 
        .A4(\read_value_mux[29][7] ), .Y(n2751) );
  OA221X1_RVT U3788 ( .A1(n1740), .A2(\read_value_mux[29][7] ), .A3(n1738), 
        .A4(\read_value_mux[29][6] ), .A5(n2751), .Y(n2758) );
  AOI22X1_RVT U3789 ( .A1(n1742), .A2(\read_value_mux[29][4] ), .A3(n1525), 
        .A4(\read_value_mux[29][5] ), .Y(n2752) );
  OA221X1_RVT U3790 ( .A1(n1745), .A2(\read_value_mux[29][5] ), .A3(n1742), 
        .A4(\read_value_mux[29][4] ), .A5(n2752), .Y(n2757) );
  AOI22X1_RVT U3791 ( .A1(n1524), .A2(\read_value_mux[29][2] ), .A3(n1750), 
        .A4(\read_value_mux[29][3] ), .Y(n2753) );
  OA221X1_RVT U3792 ( .A1(n1750), .A2(\read_value_mux[29][3] ), .A3(n1524), 
        .A4(\read_value_mux[29][2] ), .A5(n2753), .Y(n2756) );
  OA221X1_RVT U3793 ( .A1(search_data[0]), .A2(n1623), .A3(n1751), .A4(
        \read_value_mux[29][0] ), .A5(search), .Y(n2754) );
  OA221X1_RVT U3794 ( .A1(search_data[31]), .A2(n1624), .A3(n1766), .A4(
        \read_value_mux[29][31] ), .A5(n2754), .Y(n2755) );
  NAND4X0_RVT U3795 ( .A1(n2758), .A2(n2757), .A3(n2756), .A4(n2755), .Y(n2759) );
  AO22X1_RVT U3796 ( .A1(search_data[28]), .A2(\read_value_mux[31][28] ), .A3(
        n1757), .A4(n1554), .Y(n2763) );
  OA221X1_RVT U3797 ( .A1(search_data[1]), .A2(n6), .A3(n1754), .A4(
        \read_value_mux[31][1] ), .A5(n2763), .Y(n2770) );
  AO22X1_RVT U3798 ( .A1(search_data[30]), .A2(\read_value_mux[31][30] ), .A3(
        n1763), .A4(n7), .Y(n2764) );
  OA221X1_RVT U3799 ( .A1(search_data[29]), .A2(n1594), .A3(n1760), .A4(
        \read_value_mux[31][29] ), .A5(n2764), .Y(n2769) );
  AOI22X1_RVT U3800 ( .A1(n1543), .A2(\read_value_mux[31][26] ), .A3(n1542), 
        .A4(\read_value_mux[31][27] ), .Y(n2765) );
  OA221X1_RVT U3801 ( .A1(n1542), .A2(\read_value_mux[31][27] ), .A3(n1691), 
        .A4(\read_value_mux[31][26] ), .A5(n2765), .Y(n2768) );
  AOI22X1_RVT U3802 ( .A1(n1541), .A2(\read_value_mux[31][24] ), .A3(n1540), 
        .A4(\read_value_mux[31][25] ), .Y(n2766) );
  OA221X1_RVT U3803 ( .A1(n1540), .A2(\read_value_mux[31][25] ), .A3(n1695), 
        .A4(\read_value_mux[31][24] ), .A5(n2766), .Y(n2767) );
  NAND4X0_RVT U3804 ( .A1(n2770), .A2(n2769), .A3(n2768), .A4(n2767), .Y(n2798) );
  AOI22X1_RVT U3805 ( .A1(n1539), .A2(\read_value_mux[31][22] ), .A3(n1538), 
        .A4(\read_value_mux[31][23] ), .Y(n2771) );
  OA221X1_RVT U3806 ( .A1(n1538), .A2(\read_value_mux[31][23] ), .A3(n1698), 
        .A4(\read_value_mux[31][22] ), .A5(n2771), .Y(n2778) );
  AOI22X1_RVT U3807 ( .A1(n1537), .A2(\read_value_mux[31][20] ), .A3(n1536), 
        .A4(\read_value_mux[31][21] ), .Y(n2772) );
  OA221X1_RVT U3808 ( .A1(n1703), .A2(\read_value_mux[31][21] ), .A3(n1701), 
        .A4(\read_value_mux[31][20] ), .A5(n2772), .Y(n2777) );
  AOI22X1_RVT U3809 ( .A1(n1535), .A2(\read_value_mux[31][18] ), .A3(n1534), 
        .A4(\read_value_mux[31][19] ), .Y(n2773) );
  OA221X1_RVT U3810 ( .A1(n1708), .A2(\read_value_mux[31][19] ), .A3(n1705), 
        .A4(\read_value_mux[31][18] ), .A5(n2773), .Y(n2776) );
  AOI22X1_RVT U3811 ( .A1(n1533), .A2(\read_value_mux[31][16] ), .A3(n1713), 
        .A4(\read_value_mux[31][17] ), .Y(n2774) );
  OA221X1_RVT U3812 ( .A1(n1714), .A2(\read_value_mux[31][17] ), .A3(n1710), 
        .A4(\read_value_mux[31][16] ), .A5(n2774), .Y(n2775) );
  NAND4X0_RVT U3813 ( .A1(n2778), .A2(n2777), .A3(n2776), .A4(n2775), .Y(n2797) );
  AOI22X1_RVT U3814 ( .A1(n1532), .A2(\read_value_mux[31][14] ), .A3(n1720), 
        .A4(\read_value_mux[31][15] ), .Y(n2779) );
  OA221X1_RVT U3815 ( .A1(n1722), .A2(\read_value_mux[31][15] ), .A3(n1716), 
        .A4(\read_value_mux[31][14] ), .A5(n2779), .Y(n2786) );
  AOI22X1_RVT U3816 ( .A1(n1531), .A2(\read_value_mux[31][12] ), .A3(n1530), 
        .A4(\read_value_mux[31][13] ), .Y(n2780) );
  OA221X1_RVT U3817 ( .A1(n1530), .A2(\read_value_mux[31][13] ), .A3(n1724), 
        .A4(\read_value_mux[31][12] ), .A5(n2780), .Y(n2785) );
  AOI22X1_RVT U3818 ( .A1(n1529), .A2(\read_value_mux[31][10] ), .A3(n1528), 
        .A4(\read_value_mux[31][11] ), .Y(n2781) );
  OA221X1_RVT U3819 ( .A1(n1730), .A2(\read_value_mux[31][11] ), .A3(n1727), 
        .A4(\read_value_mux[31][10] ), .A5(n2781), .Y(n2784) );
  AOI22X1_RVT U3820 ( .A1(n1527), .A2(\read_value_mux[31][8] ), .A3(n1735), 
        .A4(\read_value_mux[31][9] ), .Y(n2782) );
  OA221X1_RVT U3821 ( .A1(n1736), .A2(\read_value_mux[31][9] ), .A3(n1732), 
        .A4(\read_value_mux[31][8] ), .A5(n2782), .Y(n2783) );
  NAND4X0_RVT U3822 ( .A1(n2786), .A2(n2785), .A3(n2784), .A4(n2783), .Y(n2796) );
  AOI22X1_RVT U3823 ( .A1(n1738), .A2(\read_value_mux[31][6] ), .A3(n1739), 
        .A4(\read_value_mux[31][7] ), .Y(n2787) );
  OA221X1_RVT U3824 ( .A1(n1740), .A2(\read_value_mux[31][7] ), .A3(n1738), 
        .A4(\read_value_mux[31][6] ), .A5(n2787), .Y(n2794) );
  AOI22X1_RVT U3825 ( .A1(n1526), .A2(\read_value_mux[31][4] ), .A3(n1525), 
        .A4(\read_value_mux[31][5] ), .Y(n2788) );
  OA221X1_RVT U3826 ( .A1(n1746), .A2(\read_value_mux[31][5] ), .A3(n1742), 
        .A4(\read_value_mux[31][4] ), .A5(n2788), .Y(n2793) );
  AOI22X1_RVT U3827 ( .A1(n1749), .A2(\read_value_mux[31][2] ), .A3(n1750), 
        .A4(\read_value_mux[31][3] ), .Y(n2789) );
  OA221X1_RVT U3828 ( .A1(n1750), .A2(\read_value_mux[31][3] ), .A3(n1524), 
        .A4(\read_value_mux[31][2] ), .A5(n2789), .Y(n2792) );
  OA221X1_RVT U3829 ( .A1(search_data[0]), .A2(n1595), .A3(n1751), .A4(
        \read_value_mux[31][0] ), .A5(search), .Y(n2790) );
  OA221X1_RVT U3830 ( .A1(search_data[31]), .A2(n1596), .A3(n1766), .A4(
        \read_value_mux[31][31] ), .A5(n2790), .Y(n2791) );
  NAND4X0_RVT U3831 ( .A1(n2794), .A2(n2793), .A3(n2792), .A4(n2791), .Y(n2795) );
  AO22X1_RVT U3832 ( .A1(search_data[28]), .A2(\read_value_mux[30][28] ), .A3(
        n1757), .A4(n1566), .Y(n2799) );
  OA221X1_RVT U3833 ( .A1(search_data[1]), .A2(n88), .A3(n1754), .A4(
        \read_value_mux[30][1] ), .A5(n2799), .Y(n2806) );
  AO22X1_RVT U3834 ( .A1(search_data[30]), .A2(\read_value_mux[30][30] ), .A3(
        n1763), .A4(n89), .Y(n2800) );
  OA221X1_RVT U3835 ( .A1(search_data[29]), .A2(n1625), .A3(n1760), .A4(
        \read_value_mux[30][29] ), .A5(n2800), .Y(n2805) );
  AOI22X1_RVT U3836 ( .A1(n1543), .A2(\read_value_mux[30][26] ), .A3(n1542), 
        .A4(\read_value_mux[30][27] ), .Y(n2801) );
  OA221X1_RVT U3837 ( .A1(n1542), .A2(\read_value_mux[30][27] ), .A3(n1691), 
        .A4(\read_value_mux[30][26] ), .A5(n2801), .Y(n2804) );
  AOI22X1_RVT U3838 ( .A1(n1541), .A2(\read_value_mux[30][24] ), .A3(n1540), 
        .A4(\read_value_mux[30][25] ), .Y(n2802) );
  OA221X1_RVT U3839 ( .A1(n1540), .A2(\read_value_mux[30][25] ), .A3(n1695), 
        .A4(\read_value_mux[30][24] ), .A5(n2802), .Y(n2803) );
  NAND4X0_RVT U3840 ( .A1(n2806), .A2(n2805), .A3(n2804), .A4(n2803), .Y(n2834) );
  AOI22X1_RVT U3841 ( .A1(n1539), .A2(\read_value_mux[30][22] ), .A3(n1538), 
        .A4(\read_value_mux[30][23] ), .Y(n2807) );
  OA221X1_RVT U3842 ( .A1(n1538), .A2(\read_value_mux[30][23] ), .A3(n1698), 
        .A4(\read_value_mux[30][22] ), .A5(n2807), .Y(n2814) );
  AOI22X1_RVT U3843 ( .A1(n1537), .A2(\read_value_mux[30][20] ), .A3(n1536), 
        .A4(\read_value_mux[30][21] ), .Y(n2808) );
  OA221X1_RVT U3844 ( .A1(n1703), .A2(\read_value_mux[30][21] ), .A3(n1701), 
        .A4(\read_value_mux[30][20] ), .A5(n2808), .Y(n2813) );
  AOI22X1_RVT U3845 ( .A1(n1535), .A2(\read_value_mux[30][18] ), .A3(n1534), 
        .A4(\read_value_mux[30][19] ), .Y(n2809) );
  OA221X1_RVT U3846 ( .A1(n1708), .A2(\read_value_mux[30][19] ), .A3(n1705), 
        .A4(\read_value_mux[30][18] ), .A5(n2809), .Y(n2812) );
  AOI22X1_RVT U3847 ( .A1(n1533), .A2(\read_value_mux[30][16] ), .A3(n1713), 
        .A4(\read_value_mux[30][17] ), .Y(n2810) );
  OA221X1_RVT U3848 ( .A1(n1714), .A2(\read_value_mux[30][17] ), .A3(n1710), 
        .A4(\read_value_mux[30][16] ), .A5(n2810), .Y(n2811) );
  NAND4X0_RVT U3849 ( .A1(n2814), .A2(n2813), .A3(n2812), .A4(n2811), .Y(n2833) );
  AOI22X1_RVT U3850 ( .A1(n1532), .A2(\read_value_mux[30][14] ), .A3(n1720), 
        .A4(\read_value_mux[30][15] ), .Y(n2815) );
  OA221X1_RVT U3851 ( .A1(n1722), .A2(\read_value_mux[30][15] ), .A3(n1716), 
        .A4(\read_value_mux[30][14] ), .A5(n2815), .Y(n2822) );
  AOI22X1_RVT U3852 ( .A1(n1531), .A2(\read_value_mux[30][12] ), .A3(n1530), 
        .A4(\read_value_mux[30][13] ), .Y(n2816) );
  OA221X1_RVT U3853 ( .A1(n1530), .A2(\read_value_mux[30][13] ), .A3(n1724), 
        .A4(\read_value_mux[30][12] ), .A5(n2816), .Y(n2821) );
  AOI22X1_RVT U3854 ( .A1(n1529), .A2(\read_value_mux[30][10] ), .A3(n1528), 
        .A4(\read_value_mux[30][11] ), .Y(n2817) );
  OA221X1_RVT U3855 ( .A1(n1730), .A2(\read_value_mux[30][11] ), .A3(n1727), 
        .A4(\read_value_mux[30][10] ), .A5(n2817), .Y(n2820) );
  AOI22X1_RVT U3856 ( .A1(n1527), .A2(\read_value_mux[30][8] ), .A3(n1735), 
        .A4(\read_value_mux[30][9] ), .Y(n2818) );
  OA221X1_RVT U3857 ( .A1(n1736), .A2(\read_value_mux[30][9] ), .A3(n1732), 
        .A4(\read_value_mux[30][8] ), .A5(n2818), .Y(n2819) );
  NAND4X0_RVT U3858 ( .A1(n2822), .A2(n2821), .A3(n2820), .A4(n2819), .Y(n2832) );
  AOI22X1_RVT U3859 ( .A1(n1738), .A2(\read_value_mux[30][6] ), .A3(n1739), 
        .A4(\read_value_mux[30][7] ), .Y(n2823) );
  OA221X1_RVT U3860 ( .A1(n1740), .A2(\read_value_mux[30][7] ), .A3(n1738), 
        .A4(\read_value_mux[30][6] ), .A5(n2823), .Y(n2830) );
  AOI22X1_RVT U3861 ( .A1(n1526), .A2(\read_value_mux[30][4] ), .A3(n1525), 
        .A4(\read_value_mux[30][5] ), .Y(n2824) );
  OA221X1_RVT U3862 ( .A1(n1746), .A2(\read_value_mux[30][5] ), .A3(n1742), 
        .A4(\read_value_mux[30][4] ), .A5(n2824), .Y(n2829) );
  AOI22X1_RVT U3863 ( .A1(n1524), .A2(\read_value_mux[30][2] ), .A3(n1750), 
        .A4(\read_value_mux[30][3] ), .Y(n2825) );
  OA221X1_RVT U3864 ( .A1(n1750), .A2(\read_value_mux[30][3] ), .A3(n1524), 
        .A4(\read_value_mux[30][2] ), .A5(n2825), .Y(n2828) );
  OA221X1_RVT U3865 ( .A1(search_data[0]), .A2(n1626), .A3(n1751), .A4(
        \read_value_mux[30][0] ), .A5(search), .Y(n2826) );
  OA221X1_RVT U3866 ( .A1(search_data[31]), .A2(n1674), .A3(n1766), .A4(
        \read_value_mux[30][31] ), .A5(n2826), .Y(n2827) );
  NAND4X0_RVT U3867 ( .A1(n2830), .A2(n2829), .A3(n2828), .A4(n2827), .Y(n2831) );
  OR4X1_RVT U3868 ( .A1(n2834), .A2(n2833), .A3(n2832), .A4(n2831), .Y(n2999)
         );
  AO22X1_RVT U3869 ( .A1(search_data[28]), .A2(\read_value_mux[28][28] ), .A3(
        n1757), .A4(n1555), .Y(n2835) );
  OA221X1_RVT U3870 ( .A1(search_data[1]), .A2(n83), .A3(n1754), .A4(
        \read_value_mux[28][1] ), .A5(n2835), .Y(n2842) );
  AO22X1_RVT U3871 ( .A1(search_data[30]), .A2(\read_value_mux[28][30] ), .A3(
        n1763), .A4(n84), .Y(n2836) );
  OA221X1_RVT U3872 ( .A1(search_data[29]), .A2(n1656), .A3(n1760), .A4(
        \read_value_mux[28][29] ), .A5(n2836), .Y(n2841) );
  AOI22X1_RVT U3873 ( .A1(n1543), .A2(\read_value_mux[28][26] ), .A3(n1542), 
        .A4(\read_value_mux[28][27] ), .Y(n2837) );
  OA221X1_RVT U3874 ( .A1(n1542), .A2(\read_value_mux[28][27] ), .A3(n1691), 
        .A4(\read_value_mux[28][26] ), .A5(n2837), .Y(n2840) );
  AOI22X1_RVT U3875 ( .A1(n1541), .A2(\read_value_mux[28][24] ), .A3(n1540), 
        .A4(\read_value_mux[28][25] ), .Y(n2838) );
  OA221X1_RVT U3876 ( .A1(n1540), .A2(\read_value_mux[28][25] ), .A3(n1695), 
        .A4(\read_value_mux[28][24] ), .A5(n2838), .Y(n2839) );
  NAND4X0_RVT U3877 ( .A1(n2842), .A2(n2841), .A3(n2840), .A4(n2839), .Y(n2870) );
  AOI22X1_RVT U3878 ( .A1(n1539), .A2(\read_value_mux[28][22] ), .A3(n1538), 
        .A4(\read_value_mux[28][23] ), .Y(n2843) );
  OA221X1_RVT U3879 ( .A1(n1538), .A2(\read_value_mux[28][23] ), .A3(n1698), 
        .A4(\read_value_mux[28][22] ), .A5(n2843), .Y(n2850) );
  AOI22X1_RVT U3880 ( .A1(n1537), .A2(\read_value_mux[28][20] ), .A3(n1536), 
        .A4(\read_value_mux[28][21] ), .Y(n2844) );
  OA221X1_RVT U3881 ( .A1(n1703), .A2(\read_value_mux[28][21] ), .A3(n1701), 
        .A4(\read_value_mux[28][20] ), .A5(n2844), .Y(n2849) );
  AOI22X1_RVT U3882 ( .A1(n1535), .A2(\read_value_mux[28][18] ), .A3(n1534), 
        .A4(\read_value_mux[28][19] ), .Y(n2845) );
  OA221X1_RVT U3883 ( .A1(n1708), .A2(\read_value_mux[28][19] ), .A3(n1705), 
        .A4(\read_value_mux[28][18] ), .A5(n2845), .Y(n2848) );
  AOI22X1_RVT U3884 ( .A1(n1533), .A2(\read_value_mux[28][16] ), .A3(n1713), 
        .A4(\read_value_mux[28][17] ), .Y(n2846) );
  OA221X1_RVT U3885 ( .A1(n1714), .A2(\read_value_mux[28][17] ), .A3(n1710), 
        .A4(\read_value_mux[28][16] ), .A5(n2846), .Y(n2847) );
  NAND4X0_RVT U3886 ( .A1(n2850), .A2(n2849), .A3(n2848), .A4(n2847), .Y(n2869) );
  AOI22X1_RVT U3887 ( .A1(n1532), .A2(\read_value_mux[28][14] ), .A3(n1720), 
        .A4(\read_value_mux[28][15] ), .Y(n2851) );
  OA221X1_RVT U3888 ( .A1(n1722), .A2(\read_value_mux[28][15] ), .A3(n1716), 
        .A4(\read_value_mux[28][14] ), .A5(n2851), .Y(n2858) );
  AOI22X1_RVT U3889 ( .A1(n1531), .A2(\read_value_mux[28][12] ), .A3(n1530), 
        .A4(\read_value_mux[28][13] ), .Y(n2852) );
  OA221X1_RVT U3890 ( .A1(n1530), .A2(\read_value_mux[28][13] ), .A3(n1724), 
        .A4(\read_value_mux[28][12] ), .A5(n2852), .Y(n2857) );
  AOI22X1_RVT U3891 ( .A1(n1529), .A2(\read_value_mux[28][10] ), .A3(n1528), 
        .A4(\read_value_mux[28][11] ), .Y(n2853) );
  OA221X1_RVT U3892 ( .A1(n1730), .A2(\read_value_mux[28][11] ), .A3(n1727), 
        .A4(\read_value_mux[28][10] ), .A5(n2853), .Y(n2856) );
  AOI22X1_RVT U3893 ( .A1(n1527), .A2(\read_value_mux[28][8] ), .A3(n1735), 
        .A4(\read_value_mux[28][9] ), .Y(n2854) );
  OA221X1_RVT U3894 ( .A1(n1736), .A2(\read_value_mux[28][9] ), .A3(n1732), 
        .A4(\read_value_mux[28][8] ), .A5(n2854), .Y(n2855) );
  NAND4X0_RVT U3895 ( .A1(n2858), .A2(n2857), .A3(n2856), .A4(n2855), .Y(n2868) );
  AOI22X1_RVT U3896 ( .A1(n1738), .A2(\read_value_mux[28][6] ), .A3(n1739), 
        .A4(\read_value_mux[28][7] ), .Y(n2859) );
  OA221X1_RVT U3897 ( .A1(n1740), .A2(\read_value_mux[28][7] ), .A3(n1738), 
        .A4(\read_value_mux[28][6] ), .A5(n2859), .Y(n2866) );
  AOI22X1_RVT U3898 ( .A1(n1526), .A2(\read_value_mux[28][4] ), .A3(n1525), 
        .A4(\read_value_mux[28][5] ), .Y(n2860) );
  OA221X1_RVT U3899 ( .A1(n1746), .A2(\read_value_mux[28][5] ), .A3(n1742), 
        .A4(\read_value_mux[28][4] ), .A5(n2860), .Y(n2865) );
  AOI22X1_RVT U3900 ( .A1(n1524), .A2(\read_value_mux[28][2] ), .A3(n1750), 
        .A4(\read_value_mux[28][3] ), .Y(n2861) );
  OA221X1_RVT U3901 ( .A1(n1750), .A2(\read_value_mux[28][3] ), .A3(n1524), 
        .A4(\read_value_mux[28][2] ), .A5(n2861), .Y(n2864) );
  OA221X1_RVT U3902 ( .A1(search_data[0]), .A2(n1597), .A3(n1751), .A4(
        \read_value_mux[28][0] ), .A5(search), .Y(n2862) );
  OA221X1_RVT U3903 ( .A1(search_data[31]), .A2(n1657), .A3(n1766), .A4(
        \read_value_mux[28][31] ), .A5(n2862), .Y(n2863) );
  NAND4X0_RVT U3904 ( .A1(n2866), .A2(n2865), .A3(n2864), .A4(n2863), .Y(n2867) );
  OA221X1_RVT U3905 ( .A1(n2964), .A2(n2965), .A3(n2964), .A4(n2999), .A5(
        n3002), .Y(n2907) );
  AO22X1_RVT U3906 ( .A1(search_data[28]), .A2(\read_value_mux[25][28] ), .A3(
        n1757), .A4(n1567), .Y(n2871) );
  OA221X1_RVT U3907 ( .A1(search_data[1]), .A2(n76), .A3(n1754), .A4(
        \read_value_mux[25][1] ), .A5(n2871), .Y(n2878) );
  AO22X1_RVT U3908 ( .A1(search_data[30]), .A2(\read_value_mux[25][30] ), .A3(
        n1763), .A4(n77), .Y(n2872) );
  OA221X1_RVT U3909 ( .A1(search_data[29]), .A2(n1627), .A3(n1760), .A4(
        \read_value_mux[25][29] ), .A5(n2872), .Y(n2877) );
  AOI22X1_RVT U3910 ( .A1(n1691), .A2(\read_value_mux[25][26] ), .A3(n1542), 
        .A4(\read_value_mux[25][27] ), .Y(n2873) );
  OA221X1_RVT U3911 ( .A1(n1542), .A2(\read_value_mux[25][27] ), .A3(n1691), 
        .A4(\read_value_mux[25][26] ), .A5(n2873), .Y(n2876) );
  AOI22X1_RVT U3912 ( .A1(n1695), .A2(\read_value_mux[25][24] ), .A3(n1540), 
        .A4(\read_value_mux[25][25] ), .Y(n2874) );
  OA221X1_RVT U3913 ( .A1(n1540), .A2(\read_value_mux[25][25] ), .A3(n1695), 
        .A4(\read_value_mux[25][24] ), .A5(n2874), .Y(n2875) );
  NAND4X0_RVT U3914 ( .A1(n2878), .A2(n2877), .A3(n2876), .A4(n2875), .Y(n2906) );
  AOI22X1_RVT U3915 ( .A1(n1698), .A2(\read_value_mux[25][22] ), .A3(n1538), 
        .A4(\read_value_mux[25][23] ), .Y(n2879) );
  OA221X1_RVT U3916 ( .A1(n1538), .A2(\read_value_mux[25][23] ), .A3(n1698), 
        .A4(\read_value_mux[25][22] ), .A5(n2879), .Y(n2886) );
  AOI22X1_RVT U3917 ( .A1(n1701), .A2(\read_value_mux[25][20] ), .A3(n1536), 
        .A4(\read_value_mux[25][21] ), .Y(n2880) );
  OA221X1_RVT U3918 ( .A1(n1703), .A2(\read_value_mux[25][21] ), .A3(n1701), 
        .A4(\read_value_mux[25][20] ), .A5(n2880), .Y(n2885) );
  AOI22X1_RVT U3919 ( .A1(n1705), .A2(\read_value_mux[25][18] ), .A3(n1534), 
        .A4(\read_value_mux[25][19] ), .Y(n2881) );
  OA221X1_RVT U3920 ( .A1(n1708), .A2(\read_value_mux[25][19] ), .A3(n1705), 
        .A4(\read_value_mux[25][18] ), .A5(n2881), .Y(n2884) );
  AOI22X1_RVT U3921 ( .A1(n1710), .A2(\read_value_mux[25][16] ), .A3(n1713), 
        .A4(\read_value_mux[25][17] ), .Y(n2882) );
  OA221X1_RVT U3922 ( .A1(n1714), .A2(\read_value_mux[25][17] ), .A3(n1710), 
        .A4(\read_value_mux[25][16] ), .A5(n2882), .Y(n2883) );
  NAND4X0_RVT U3923 ( .A1(n2886), .A2(n2885), .A3(n2884), .A4(n2883), .Y(n2905) );
  AOI22X1_RVT U3924 ( .A1(n1716), .A2(\read_value_mux[25][14] ), .A3(n1720), 
        .A4(\read_value_mux[25][15] ), .Y(n2887) );
  OA221X1_RVT U3925 ( .A1(n1722), .A2(\read_value_mux[25][15] ), .A3(n1716), 
        .A4(\read_value_mux[25][14] ), .A5(n2887), .Y(n2894) );
  AOI22X1_RVT U3926 ( .A1(n1724), .A2(\read_value_mux[25][12] ), .A3(n1530), 
        .A4(\read_value_mux[25][13] ), .Y(n2888) );
  OA221X1_RVT U3927 ( .A1(n1530), .A2(\read_value_mux[25][13] ), .A3(n1724), 
        .A4(\read_value_mux[25][12] ), .A5(n2888), .Y(n2893) );
  AOI22X1_RVT U3928 ( .A1(n1727), .A2(\read_value_mux[25][10] ), .A3(n1528), 
        .A4(\read_value_mux[25][11] ), .Y(n2889) );
  OA221X1_RVT U3929 ( .A1(n1730), .A2(\read_value_mux[25][11] ), .A3(n1727), 
        .A4(\read_value_mux[25][10] ), .A5(n2889), .Y(n2892) );
  AOI22X1_RVT U3930 ( .A1(n1732), .A2(\read_value_mux[25][8] ), .A3(n1735), 
        .A4(\read_value_mux[25][9] ), .Y(n2890) );
  OA221X1_RVT U3931 ( .A1(n1736), .A2(\read_value_mux[25][9] ), .A3(n1732), 
        .A4(\read_value_mux[25][8] ), .A5(n2890), .Y(n2891) );
  NAND4X0_RVT U3932 ( .A1(n2894), .A2(n2893), .A3(n2892), .A4(n2891), .Y(n2904) );
  AOI22X1_RVT U3933 ( .A1(n2940), .A2(\read_value_mux[25][6] ), .A3(n1739), 
        .A4(\read_value_mux[25][7] ), .Y(n2895) );
  OA221X1_RVT U3934 ( .A1(n1740), .A2(\read_value_mux[25][7] ), .A3(n1738), 
        .A4(\read_value_mux[25][6] ), .A5(n2895), .Y(n2902) );
  AOI22X1_RVT U3935 ( .A1(n1742), .A2(\read_value_mux[25][4] ), .A3(n1525), 
        .A4(\read_value_mux[25][5] ), .Y(n2896) );
  OA221X1_RVT U3936 ( .A1(n1746), .A2(\read_value_mux[25][5] ), .A3(n1742), 
        .A4(\read_value_mux[25][4] ), .A5(n2896), .Y(n2901) );
  AOI22X1_RVT U3937 ( .A1(n1524), .A2(\read_value_mux[25][2] ), .A3(n1750), 
        .A4(\read_value_mux[25][3] ), .Y(n2897) );
  OA221X1_RVT U3938 ( .A1(n1750), .A2(\read_value_mux[25][3] ), .A3(n1524), 
        .A4(\read_value_mux[25][2] ), .A5(n2897), .Y(n2900) );
  OA221X1_RVT U3939 ( .A1(search_data[0]), .A2(n1628), .A3(n1751), .A4(
        \read_value_mux[25][0] ), .A5(search), .Y(n2898) );
  OA221X1_RVT U3940 ( .A1(search_data[31]), .A2(n1629), .A3(n1766), .A4(
        \read_value_mux[25][31] ), .A5(n2898), .Y(n2899) );
  NAND4X0_RVT U3941 ( .A1(n2902), .A2(n2901), .A3(n2900), .A4(n2899), .Y(n2903) );
  AO22X1_RVT U3942 ( .A1(search_data[28]), .A2(\read_value_mux[8][28] ), .A3(
        n1758), .A4(n1556), .Y(n2908) );
  OA221X1_RVT U3943 ( .A1(search_data[1]), .A2(n30), .A3(n1755), .A4(
        \read_value_mux[8][1] ), .A5(n2908), .Y(n2916) );
  AO22X1_RVT U3944 ( .A1(search_data[30]), .A2(\read_value_mux[8][30] ), .A3(
        n1764), .A4(n31), .Y(n2909) );
  OA221X1_RVT U3945 ( .A1(search_data[29]), .A2(n1598), .A3(n1761), .A4(
        \read_value_mux[8][29] ), .A5(n2909), .Y(n2915) );
  AOI22X1_RVT U3946 ( .A1(n1543), .A2(\read_value_mux[8][26] ), .A3(n1542), 
        .A4(\read_value_mux[8][27] ), .Y(n2910) );
  OA221X1_RVT U3947 ( .A1(n1542), .A2(\read_value_mux[8][27] ), .A3(n1691), 
        .A4(\read_value_mux[8][26] ), .A5(n2910), .Y(n2914) );
  AOI22X1_RVT U3948 ( .A1(n1541), .A2(\read_value_mux[8][24] ), .A3(n1540), 
        .A4(\read_value_mux[8][25] ), .Y(n2911) );
  OA221X1_RVT U3949 ( .A1(n1697), .A2(\read_value_mux[8][25] ), .A3(n1695), 
        .A4(\read_value_mux[8][24] ), .A5(n2911), .Y(n2913) );
  NAND4X0_RVT U3950 ( .A1(n2916), .A2(n2915), .A3(n2914), .A4(n2913), .Y(n2952) );
  AOI22X1_RVT U3951 ( .A1(n1539), .A2(\read_value_mux[8][22] ), .A3(n1538), 
        .A4(\read_value_mux[8][23] ), .Y(n2917) );
  OA221X1_RVT U3952 ( .A1(n1538), .A2(\read_value_mux[8][23] ), .A3(n1698), 
        .A4(\read_value_mux[8][22] ), .A5(n2917), .Y(n2927) );
  AOI22X1_RVT U3953 ( .A1(n1537), .A2(\read_value_mux[8][20] ), .A3(n1536), 
        .A4(\read_value_mux[8][21] ), .Y(n2919) );
  OA221X1_RVT U3954 ( .A1(n1704), .A2(\read_value_mux[8][21] ), .A3(n1701), 
        .A4(\read_value_mux[8][20] ), .A5(n2919), .Y(n2926) );
  AOI22X1_RVT U3955 ( .A1(n1535), .A2(\read_value_mux[8][18] ), .A3(n1534), 
        .A4(\read_value_mux[8][19] ), .Y(n2921) );
  OA221X1_RVT U3956 ( .A1(n1709), .A2(\read_value_mux[8][19] ), .A3(n1705), 
        .A4(\read_value_mux[8][18] ), .A5(n2921), .Y(n2925) );
  AOI22X1_RVT U3957 ( .A1(n1533), .A2(\read_value_mux[8][16] ), .A3(n1713), 
        .A4(\read_value_mux[8][17] ), .Y(n2922) );
  OA221X1_RVT U3958 ( .A1(n1715), .A2(\read_value_mux[8][17] ), .A3(n1710), 
        .A4(\read_value_mux[8][16] ), .A5(n2922), .Y(n2924) );
  NAND4X0_RVT U3959 ( .A1(n2927), .A2(n2926), .A3(n2925), .A4(n2924), .Y(n2951) );
  AOI22X1_RVT U3960 ( .A1(n1532), .A2(\read_value_mux[8][14] ), .A3(n1720), 
        .A4(\read_value_mux[8][15] ), .Y(n2928) );
  OA221X1_RVT U3961 ( .A1(n1723), .A2(\read_value_mux[8][15] ), .A3(n1716), 
        .A4(\read_value_mux[8][14] ), .A5(n2928), .Y(n2938) );
  AOI22X1_RVT U3962 ( .A1(n1531), .A2(\read_value_mux[8][12] ), .A3(n1530), 
        .A4(\read_value_mux[8][13] ), .Y(n2930) );
  OA221X1_RVT U3963 ( .A1(n1530), .A2(\read_value_mux[8][13] ), .A3(n1724), 
        .A4(\read_value_mux[8][12] ), .A5(n2930), .Y(n2937) );
  AOI22X1_RVT U3964 ( .A1(n1529), .A2(\read_value_mux[8][10] ), .A3(n1528), 
        .A4(\read_value_mux[8][11] ), .Y(n2932) );
  OA221X1_RVT U3965 ( .A1(n1731), .A2(\read_value_mux[8][11] ), .A3(n1727), 
        .A4(\read_value_mux[8][10] ), .A5(n2932), .Y(n2936) );
  AOI22X1_RVT U3966 ( .A1(n1527), .A2(\read_value_mux[8][8] ), .A3(n1735), 
        .A4(\read_value_mux[8][9] ), .Y(n2933) );
  OA221X1_RVT U3967 ( .A1(n1737), .A2(\read_value_mux[8][9] ), .A3(n1732), 
        .A4(\read_value_mux[8][8] ), .A5(n2933), .Y(n2935) );
  NAND4X0_RVT U3968 ( .A1(n2938), .A2(n2937), .A3(n2936), .A4(n2935), .Y(n2950) );
  AOI22X1_RVT U3969 ( .A1(n2940), .A2(\read_value_mux[8][6] ), .A3(n1739), 
        .A4(\read_value_mux[8][7] ), .Y(n2939) );
  OA221X1_RVT U3970 ( .A1(n1741), .A2(\read_value_mux[8][7] ), .A3(n1738), 
        .A4(\read_value_mux[8][6] ), .A5(n2939), .Y(n2948) );
  AOI22X1_RVT U3971 ( .A1(n1526), .A2(\read_value_mux[8][4] ), .A3(n1525), 
        .A4(\read_value_mux[8][5] ), .Y(n2941) );
  OA221X1_RVT U3972 ( .A1(n1747), .A2(\read_value_mux[8][5] ), .A3(n1742), 
        .A4(\read_value_mux[8][4] ), .A5(n2941), .Y(n2947) );
  AOI22X1_RVT U3973 ( .A1(n1524), .A2(\read_value_mux[8][2] ), .A3(n1750), 
        .A4(\read_value_mux[8][3] ), .Y(n2943) );
  OA221X1_RVT U3974 ( .A1(n1750), .A2(\read_value_mux[8][3] ), .A3(n1524), 
        .A4(\read_value_mux[8][2] ), .A5(n2943), .Y(n2946) );
  OA221X1_RVT U3975 ( .A1(search_data[0]), .A2(n1599), .A3(n1752), .A4(
        \read_value_mux[8][0] ), .A5(search), .Y(n2944) );
  OA221X1_RVT U3976 ( .A1(search_data[31]), .A2(n1600), .A3(n1767), .A4(
        \read_value_mux[8][31] ), .A5(n2944), .Y(n2945) );
  NAND4X0_RVT U3977 ( .A1(n2948), .A2(n2947), .A3(n2946), .A4(n2945), .Y(n2949) );
  NAND2X0_RVT U3978 ( .A1(n3012), .A2(n3011), .Y(n2953) );
  NAND2X0_RVT U3979 ( .A1(n2994), .A2(n2993), .Y(n3105) );
  NAND2X0_RVT U3980 ( .A1(n3000), .A2(n2999), .Y(n2966) );
  NAND4X0_RVT U3981 ( .A1(n3101), .A2(n3002), .A3(n3001), .A4(n2966), .Y(n2967) );
  NAND3X0_RVT U3982 ( .A1(n3103), .A2(n3102), .A3(n2967), .Y(n2968) );
  AND4X1_RVT U3983 ( .A1(n3104), .A2(n2985), .A3(n2996), .A4(n2968), .Y(n2972)
         );
  NAND2X0_RVT U3984 ( .A1(n2971), .A2(n2970), .Y(n3107) );
  AND2X1_RVT U3985 ( .A1(n2975), .A2(n2974), .Y(n2991) );
  NAND2X0_RVT U3986 ( .A1(n3100), .A2(n3099), .Y(n2981) );
  NAND3X0_RVT U3987 ( .A1(n3101), .A2(n3104), .A3(n2981), .Y(n2982) );
  NAND3X0_RVT U3988 ( .A1(n2983), .A2(n2997), .A3(n2982), .Y(n2984) );
  AND2X1_RVT U3989 ( .A1(n2992), .A2(n2991), .Y(n3109) );
  NAND4X0_RVT U3990 ( .A1(n2995), .A2(n3109), .A3(n2994), .A4(n2993), .Y(n3014) );
  AND3X1_RVT U3991 ( .A1(n2998), .A2(n2997), .A3(n2996), .Y(n3106) );
  NAND4X0_RVT U3992 ( .A1(n3002), .A2(n3001), .A3(n3000), .A4(n2999), .Y(n3098) );
  NAND4X0_RVT U3993 ( .A1(n3101), .A2(n3003), .A3(n3100), .A4(n3099), .Y(n3015) );
  NAND4X0_RVT U3994 ( .A1(n3012), .A2(n3011), .A3(n3010), .A4(n3009), .Y(n3110) );
  AO22X1_RVT U3995 ( .A1(\read_value_mux[0][0] ), .A2(n1675), .A3(
        write_data[0]), .A4(n3019), .Y(\words[0]/data_i[0] ) );
  AO22X1_RVT U3996 ( .A1(\read_value_mux[0][10] ), .A2(n1675), .A3(n3019), 
        .A4(write_data[10]), .Y(\words[0]/data_i[10] ) );
  AO22X1_RVT U3997 ( .A1(\read_value_mux[0][11] ), .A2(n1675), .A3(n3019), 
        .A4(write_data[11]), .Y(\words[0]/data_i[11] ) );
  AO22X1_RVT U3998 ( .A1(\read_value_mux[0][12] ), .A2(n1675), .A3(n3019), 
        .A4(write_data[12]), .Y(\words[0]/data_i[12] ) );
  AO22X1_RVT U3999 ( .A1(\read_value_mux[0][13] ), .A2(n1675), .A3(n3019), 
        .A4(write_data[13]), .Y(\words[0]/data_i[13] ) );
  AO22X1_RVT U4000 ( .A1(\read_value_mux[0][14] ), .A2(n1675), .A3(n3019), 
        .A4(write_data[14]), .Y(\words[0]/data_i[14] ) );
  AO22X1_RVT U4001 ( .A1(\read_value_mux[0][15] ), .A2(n1675), .A3(n3019), 
        .A4(write_data[15]), .Y(\words[0]/data_i[15] ) );
  AO22X1_RVT U4002 ( .A1(\read_value_mux[0][16] ), .A2(n1675), .A3(n3019), 
        .A4(write_data[16]), .Y(\words[0]/data_i[16] ) );
  AO22X1_RVT U4003 ( .A1(\read_value_mux[0][17] ), .A2(n1675), .A3(n3019), 
        .A4(write_data[17]), .Y(\words[0]/data_i[17] ) );
  AO22X1_RVT U4004 ( .A1(\read_value_mux[0][18] ), .A2(n1675), .A3(n3019), 
        .A4(write_data[18]), .Y(\words[0]/data_i[18] ) );
  AO22X1_RVT U4005 ( .A1(\read_value_mux[0][19] ), .A2(n1675), .A3(n3019), 
        .A4(write_data[19]), .Y(\words[0]/data_i[19] ) );
  AO22X1_RVT U4006 ( .A1(write_data[1]), .A2(n3019), .A3(
        \read_value_mux[0][1] ), .A4(n1675), .Y(\words[0]/data_i[1] ) );
  AO22X1_RVT U4007 ( .A1(\read_value_mux[0][20] ), .A2(n1675), .A3(n3019), 
        .A4(write_data[20]), .Y(\words[0]/data_i[20] ) );
  AO22X1_RVT U4008 ( .A1(\read_value_mux[0][21] ), .A2(n1675), .A3(n3019), 
        .A4(write_data[21]), .Y(\words[0]/data_i[21] ) );
  AO22X1_RVT U4009 ( .A1(\read_value_mux[0][22] ), .A2(n1675), .A3(n3019), 
        .A4(write_data[22]), .Y(\words[0]/data_i[22] ) );
  AO22X1_RVT U4010 ( .A1(\read_value_mux[0][23] ), .A2(n1675), .A3(n3019), 
        .A4(write_data[23]), .Y(\words[0]/data_i[23] ) );
  AO22X1_RVT U4011 ( .A1(\read_value_mux[0][24] ), .A2(n1675), .A3(n3019), 
        .A4(write_data[24]), .Y(\words[0]/data_i[24] ) );
  AO22X1_RVT U4012 ( .A1(\read_value_mux[0][25] ), .A2(n1675), .A3(n3019), 
        .A4(write_data[25]), .Y(\words[0]/data_i[25] ) );
  AO22X1_RVT U4013 ( .A1(\read_value_mux[0][26] ), .A2(n1675), .A3(n3019), 
        .A4(write_data[26]), .Y(\words[0]/data_i[26] ) );
  AO22X1_RVT U4014 ( .A1(\read_value_mux[0][27] ), .A2(n1675), .A3(n3019), 
        .A4(write_data[27]), .Y(\words[0]/data_i[27] ) );
  AO22X1_RVT U4015 ( .A1(\read_value_mux[0][28] ), .A2(n1675), .A3(n3019), 
        .A4(write_data[28]), .Y(\words[0]/data_i[28] ) );
  AO22X1_RVT U4016 ( .A1(\read_value_mux[0][29] ), .A2(n1675), .A3(n3019), 
        .A4(write_data[29]), .Y(\words[0]/data_i[29] ) );
  AO22X1_RVT U4017 ( .A1(\read_value_mux[0][2] ), .A2(n1675), .A3(n3019), .A4(
        write_data[2]), .Y(\words[0]/data_i[2] ) );
  AO22X1_RVT U4018 ( .A1(write_data[30]), .A2(n3019), .A3(
        \read_value_mux[0][30] ), .A4(n1675), .Y(\words[0]/data_i[30] ) );
  AO22X1_RVT U4019 ( .A1(\read_value_mux[0][31] ), .A2(n1675), .A3(n3019), 
        .A4(write_data[31]), .Y(\words[0]/data_i[31] ) );
  AO22X1_RVT U4020 ( .A1(\read_value_mux[0][3] ), .A2(n1675), .A3(n3019), .A4(
        write_data[3]), .Y(\words[0]/data_i[3] ) );
  AO22X1_RVT U4021 ( .A1(\read_value_mux[0][4] ), .A2(n1675), .A3(n3019), .A4(
        write_data[4]), .Y(\words[0]/data_i[4] ) );
  AO22X1_RVT U4022 ( .A1(\read_value_mux[0][5] ), .A2(n1675), .A3(n3019), .A4(
        write_data[5]), .Y(\words[0]/data_i[5] ) );
  AO22X1_RVT U4023 ( .A1(\read_value_mux[0][6] ), .A2(n1675), .A3(n3019), .A4(
        write_data[6]), .Y(\words[0]/data_i[6] ) );
  AO22X1_RVT U4024 ( .A1(\read_value_mux[0][7] ), .A2(n1675), .A3(n3019), .A4(
        write_data[7]), .Y(\words[0]/data_i[7] ) );
  AO22X1_RVT U4025 ( .A1(\read_value_mux[0][8] ), .A2(n1675), .A3(n3019), .A4(
        write_data[8]), .Y(\words[0]/data_i[8] ) );
  AO22X1_RVT U4026 ( .A1(\read_value_mux[0][9] ), .A2(n1675), .A3(n3019), .A4(
        write_data[9]), .Y(\words[0]/data_i[9] ) );
  AO21X1_RVT U4027 ( .A1(\words[0]/valid_o ), .A2(n1675), .A3(n3019), .Y(
        \words[0]/valid_i ) );
  AO22X1_RVT U4028 ( .A1(\read_value_mux[10][0] ), .A2(n1685), .A3(
        write_data[0]), .A4(n3021), .Y(\words[10]/data_i[0] ) );
  AO22X1_RVT U4029 ( .A1(\read_value_mux[10][10] ), .A2(n1685), .A3(
        write_data[10]), .A4(n3021), .Y(\words[10]/data_i[10] ) );
  AO22X1_RVT U4030 ( .A1(\read_value_mux[10][11] ), .A2(n1685), .A3(
        write_data[11]), .A4(n3021), .Y(\words[10]/data_i[11] ) );
  AO22X1_RVT U4031 ( .A1(\read_value_mux[10][12] ), .A2(n1685), .A3(
        write_data[12]), .A4(n3021), .Y(\words[10]/data_i[12] ) );
  AO22X1_RVT U4032 ( .A1(\read_value_mux[10][13] ), .A2(n1685), .A3(
        write_data[13]), .A4(n3021), .Y(\words[10]/data_i[13] ) );
  AO22X1_RVT U4033 ( .A1(\read_value_mux[10][14] ), .A2(n1685), .A3(
        write_data[14]), .A4(n3021), .Y(\words[10]/data_i[14] ) );
  AO22X1_RVT U4034 ( .A1(\read_value_mux[10][15] ), .A2(n1685), .A3(
        write_data[15]), .A4(n3021), .Y(\words[10]/data_i[15] ) );
  AO22X1_RVT U4035 ( .A1(\read_value_mux[10][16] ), .A2(n1685), .A3(
        write_data[16]), .A4(n3021), .Y(\words[10]/data_i[16] ) );
  AO22X1_RVT U4036 ( .A1(\read_value_mux[10][17] ), .A2(n1685), .A3(
        write_data[17]), .A4(n3021), .Y(\words[10]/data_i[17] ) );
  AO22X1_RVT U4037 ( .A1(\read_value_mux[10][18] ), .A2(n1685), .A3(
        write_data[18]), .A4(n3021), .Y(\words[10]/data_i[18] ) );
  AO22X1_RVT U4038 ( .A1(\read_value_mux[10][19] ), .A2(n1685), .A3(
        write_data[19]), .A4(n3021), .Y(\words[10]/data_i[19] ) );
  AO22X1_RVT U4039 ( .A1(n3021), .A2(write_data[1]), .A3(
        \read_value_mux[10][1] ), .A4(n1685), .Y(\words[10]/data_i[1] ) );
  AO22X1_RVT U4040 ( .A1(\read_value_mux[10][20] ), .A2(n1685), .A3(
        write_data[20]), .A4(n3021), .Y(\words[10]/data_i[20] ) );
  AO22X1_RVT U4041 ( .A1(\read_value_mux[10][21] ), .A2(n1685), .A3(
        write_data[21]), .A4(n3021), .Y(\words[10]/data_i[21] ) );
  AO22X1_RVT U4042 ( .A1(\read_value_mux[10][22] ), .A2(n1685), .A3(
        write_data[22]), .A4(n3021), .Y(\words[10]/data_i[22] ) );
  AO22X1_RVT U4043 ( .A1(\read_value_mux[10][23] ), .A2(n1685), .A3(
        write_data[23]), .A4(n3021), .Y(\words[10]/data_i[23] ) );
  AO22X1_RVT U4044 ( .A1(\read_value_mux[10][24] ), .A2(n1685), .A3(
        write_data[24]), .A4(n3021), .Y(\words[10]/data_i[24] ) );
  AO22X1_RVT U4045 ( .A1(\read_value_mux[10][25] ), .A2(n1685), .A3(
        write_data[25]), .A4(n3021), .Y(\words[10]/data_i[25] ) );
  AO22X1_RVT U4046 ( .A1(\read_value_mux[10][26] ), .A2(n1685), .A3(
        write_data[26]), .A4(n3021), .Y(\words[10]/data_i[26] ) );
  AO22X1_RVT U4047 ( .A1(\read_value_mux[10][27] ), .A2(n1685), .A3(
        write_data[27]), .A4(n3021), .Y(\words[10]/data_i[27] ) );
  AO22X1_RVT U4048 ( .A1(\read_value_mux[10][28] ), .A2(n1685), .A3(
        write_data[28]), .A4(n3021), .Y(\words[10]/data_i[28] ) );
  AO22X1_RVT U4049 ( .A1(\read_value_mux[10][29] ), .A2(n1685), .A3(
        write_data[29]), .A4(n3021), .Y(\words[10]/data_i[29] ) );
  AO22X1_RVT U4050 ( .A1(\read_value_mux[10][2] ), .A2(n1685), .A3(
        write_data[2]), .A4(n3021), .Y(\words[10]/data_i[2] ) );
  AO22X1_RVT U4051 ( .A1(n3021), .A2(write_data[30]), .A3(
        \read_value_mux[10][30] ), .A4(n1685), .Y(\words[10]/data_i[30] ) );
  AO22X1_RVT U4052 ( .A1(\read_value_mux[10][31] ), .A2(n1685), .A3(
        write_data[31]), .A4(n3021), .Y(\words[10]/data_i[31] ) );
  AO22X1_RVT U4053 ( .A1(\read_value_mux[10][3] ), .A2(n1685), .A3(
        write_data[3]), .A4(n3021), .Y(\words[10]/data_i[3] ) );
  AO22X1_RVT U4054 ( .A1(\read_value_mux[10][4] ), .A2(n1685), .A3(
        write_data[4]), .A4(n3021), .Y(\words[10]/data_i[4] ) );
  AO22X1_RVT U4055 ( .A1(\read_value_mux[10][5] ), .A2(n1685), .A3(
        write_data[5]), .A4(n3021), .Y(\words[10]/data_i[5] ) );
  AO22X1_RVT U4056 ( .A1(\read_value_mux[10][6] ), .A2(n1685), .A3(
        write_data[6]), .A4(n3021), .Y(\words[10]/data_i[6] ) );
  AO22X1_RVT U4057 ( .A1(\read_value_mux[10][7] ), .A2(n1685), .A3(
        write_data[7]), .A4(n3021), .Y(\words[10]/data_i[7] ) );
  AO22X1_RVT U4058 ( .A1(\read_value_mux[10][8] ), .A2(n1685), .A3(
        write_data[8]), .A4(n3021), .Y(\words[10]/data_i[8] ) );
  AO22X1_RVT U4059 ( .A1(\read_value_mux[10][9] ), .A2(n1685), .A3(
        write_data[9]), .A4(n3021), .Y(\words[10]/data_i[9] ) );
  AO21X1_RVT U4060 ( .A1(\words[10]/valid_o ), .A2(n1685), .A3(n3021), .Y(
        \words[10]/valid_i ) );
  AO22X1_RVT U4061 ( .A1(\read_value_mux[11][0] ), .A2(n1686), .A3(
        write_data[0]), .A4(n3023), .Y(\words[11]/data_i[0] ) );
  AO22X1_RVT U4062 ( .A1(\read_value_mux[11][10] ), .A2(n1686), .A3(
        write_data[10]), .A4(n3023), .Y(\words[11]/data_i[10] ) );
  AO22X1_RVT U4063 ( .A1(\read_value_mux[11][11] ), .A2(n1686), .A3(
        write_data[11]), .A4(n3023), .Y(\words[11]/data_i[11] ) );
  AO22X1_RVT U4064 ( .A1(\read_value_mux[11][12] ), .A2(n1686), .A3(
        write_data[12]), .A4(n3023), .Y(\words[11]/data_i[12] ) );
  AO22X1_RVT U4065 ( .A1(\read_value_mux[11][13] ), .A2(n1686), .A3(
        write_data[13]), .A4(n3023), .Y(\words[11]/data_i[13] ) );
  AO22X1_RVT U4066 ( .A1(\read_value_mux[11][14] ), .A2(n1686), .A3(
        write_data[14]), .A4(n3023), .Y(\words[11]/data_i[14] ) );
  AO22X1_RVT U4067 ( .A1(\read_value_mux[11][15] ), .A2(n1686), .A3(
        write_data[15]), .A4(n3023), .Y(\words[11]/data_i[15] ) );
  AO22X1_RVT U4068 ( .A1(\read_value_mux[11][16] ), .A2(n1686), .A3(
        write_data[16]), .A4(n3023), .Y(\words[11]/data_i[16] ) );
  AO22X1_RVT U4069 ( .A1(\read_value_mux[11][17] ), .A2(n1686), .A3(
        write_data[17]), .A4(n3023), .Y(\words[11]/data_i[17] ) );
  AO22X1_RVT U4070 ( .A1(\read_value_mux[11][18] ), .A2(n1686), .A3(
        write_data[18]), .A4(n3023), .Y(\words[11]/data_i[18] ) );
  AO22X1_RVT U4071 ( .A1(\read_value_mux[11][19] ), .A2(n1686), .A3(
        write_data[19]), .A4(n3023), .Y(\words[11]/data_i[19] ) );
  AO22X1_RVT U4072 ( .A1(n3023), .A2(write_data[1]), .A3(
        \read_value_mux[11][1] ), .A4(n1686), .Y(\words[11]/data_i[1] ) );
  AO22X1_RVT U4073 ( .A1(\read_value_mux[11][20] ), .A2(n1686), .A3(
        write_data[20]), .A4(n3023), .Y(\words[11]/data_i[20] ) );
  AO22X1_RVT U4074 ( .A1(\read_value_mux[11][21] ), .A2(n1686), .A3(
        write_data[21]), .A4(n3023), .Y(\words[11]/data_i[21] ) );
  AO22X1_RVT U4075 ( .A1(\read_value_mux[11][22] ), .A2(n1686), .A3(
        write_data[22]), .A4(n3023), .Y(\words[11]/data_i[22] ) );
  AO22X1_RVT U4076 ( .A1(\read_value_mux[11][23] ), .A2(n1686), .A3(
        write_data[23]), .A4(n3023), .Y(\words[11]/data_i[23] ) );
  AO22X1_RVT U4077 ( .A1(\read_value_mux[11][24] ), .A2(n1686), .A3(
        write_data[24]), .A4(n3023), .Y(\words[11]/data_i[24] ) );
  AO22X1_RVT U4078 ( .A1(\read_value_mux[11][25] ), .A2(n1686), .A3(
        write_data[25]), .A4(n3023), .Y(\words[11]/data_i[25] ) );
  AO22X1_RVT U4079 ( .A1(\read_value_mux[11][26] ), .A2(n1686), .A3(
        write_data[26]), .A4(n3023), .Y(\words[11]/data_i[26] ) );
  AO22X1_RVT U4080 ( .A1(\read_value_mux[11][27] ), .A2(n1686), .A3(
        write_data[27]), .A4(n3023), .Y(\words[11]/data_i[27] ) );
  AO22X1_RVT U4081 ( .A1(\read_value_mux[11][28] ), .A2(n1686), .A3(
        write_data[28]), .A4(n3023), .Y(\words[11]/data_i[28] ) );
  AO22X1_RVT U4082 ( .A1(\read_value_mux[11][29] ), .A2(n1686), .A3(
        write_data[29]), .A4(n3023), .Y(\words[11]/data_i[29] ) );
  AO22X1_RVT U4083 ( .A1(\read_value_mux[11][2] ), .A2(n1686), .A3(
        write_data[2]), .A4(n3023), .Y(\words[11]/data_i[2] ) );
  AO22X1_RVT U4084 ( .A1(n3023), .A2(write_data[30]), .A3(
        \read_value_mux[11][30] ), .A4(n1686), .Y(\words[11]/data_i[30] ) );
  AO22X1_RVT U4085 ( .A1(\read_value_mux[11][31] ), .A2(n1686), .A3(
        write_data[31]), .A4(n3023), .Y(\words[11]/data_i[31] ) );
  AO22X1_RVT U4086 ( .A1(\read_value_mux[11][3] ), .A2(n1686), .A3(
        write_data[3]), .A4(n3023), .Y(\words[11]/data_i[3] ) );
  AO22X1_RVT U4087 ( .A1(\read_value_mux[11][4] ), .A2(n1686), .A3(
        write_data[4]), .A4(n3023), .Y(\words[11]/data_i[4] ) );
  AO22X1_RVT U4088 ( .A1(\read_value_mux[11][5] ), .A2(n1686), .A3(
        write_data[5]), .A4(n3023), .Y(\words[11]/data_i[5] ) );
  AO22X1_RVT U4089 ( .A1(\read_value_mux[11][6] ), .A2(n1686), .A3(
        write_data[6]), .A4(n3023), .Y(\words[11]/data_i[6] ) );
  AO22X1_RVT U4090 ( .A1(\read_value_mux[11][7] ), .A2(n1686), .A3(
        write_data[7]), .A4(n3023), .Y(\words[11]/data_i[7] ) );
  AO22X1_RVT U4091 ( .A1(\read_value_mux[11][8] ), .A2(n1686), .A3(
        write_data[8]), .A4(n3023), .Y(\words[11]/data_i[8] ) );
  AO22X1_RVT U4092 ( .A1(\read_value_mux[11][9] ), .A2(n1686), .A3(
        write_data[9]), .A4(n3023), .Y(\words[11]/data_i[9] ) );
  AO21X1_RVT U4093 ( .A1(\words[11]/valid_o ), .A2(n1686), .A3(n3023), .Y(
        \words[11]/valid_i ) );
  AO22X1_RVT U4094 ( .A1(\read_value_mux[12][0] ), .A2(n3025), .A3(
        write_data[0]), .A4(n3024), .Y(\words[12]/data_i[0] ) );
  AO22X1_RVT U4095 ( .A1(\read_value_mux[12][10] ), .A2(n3025), .A3(
        write_data[10]), .A4(n3024), .Y(\words[12]/data_i[10] ) );
  AO22X1_RVT U4096 ( .A1(\read_value_mux[12][11] ), .A2(n3025), .A3(
        write_data[11]), .A4(n3024), .Y(\words[12]/data_i[11] ) );
  AO22X1_RVT U4097 ( .A1(\read_value_mux[12][12] ), .A2(n3025), .A3(
        write_data[12]), .A4(n3024), .Y(\words[12]/data_i[12] ) );
  AO22X1_RVT U4098 ( .A1(\read_value_mux[12][13] ), .A2(n3025), .A3(
        write_data[13]), .A4(n3024), .Y(\words[12]/data_i[13] ) );
  AO22X1_RVT U4099 ( .A1(\read_value_mux[12][14] ), .A2(n3025), .A3(
        write_data[14]), .A4(n3024), .Y(\words[12]/data_i[14] ) );
  AO22X1_RVT U4100 ( .A1(\read_value_mux[12][15] ), .A2(n3025), .A3(
        write_data[15]), .A4(n3024), .Y(\words[12]/data_i[15] ) );
  AO22X1_RVT U4101 ( .A1(\read_value_mux[12][16] ), .A2(n3025), .A3(
        write_data[16]), .A4(n3024), .Y(\words[12]/data_i[16] ) );
  AO22X1_RVT U4102 ( .A1(\read_value_mux[12][17] ), .A2(n3025), .A3(
        write_data[17]), .A4(n3024), .Y(\words[12]/data_i[17] ) );
  AO22X1_RVT U4103 ( .A1(\read_value_mux[12][18] ), .A2(n3025), .A3(
        write_data[18]), .A4(n3024), .Y(\words[12]/data_i[18] ) );
  AO22X1_RVT U4104 ( .A1(\read_value_mux[12][19] ), .A2(n3025), .A3(
        write_data[19]), .A4(n3024), .Y(\words[12]/data_i[19] ) );
  AO22X1_RVT U4105 ( .A1(n3024), .A2(write_data[1]), .A3(
        \read_value_mux[12][1] ), .A4(n3025), .Y(\words[12]/data_i[1] ) );
  AO22X1_RVT U4106 ( .A1(\read_value_mux[12][20] ), .A2(n3025), .A3(
        write_data[20]), .A4(n3024), .Y(\words[12]/data_i[20] ) );
  AO22X1_RVT U4107 ( .A1(\read_value_mux[12][21] ), .A2(n3025), .A3(
        write_data[21]), .A4(n3024), .Y(\words[12]/data_i[21] ) );
  AO22X1_RVT U4108 ( .A1(\read_value_mux[12][22] ), .A2(n3025), .A3(
        write_data[22]), .A4(n3024), .Y(\words[12]/data_i[22] ) );
  AO22X1_RVT U4109 ( .A1(\read_value_mux[12][23] ), .A2(n3025), .A3(
        write_data[23]), .A4(n3024), .Y(\words[12]/data_i[23] ) );
  AO22X1_RVT U4110 ( .A1(\read_value_mux[12][24] ), .A2(n3025), .A3(
        write_data[24]), .A4(n3024), .Y(\words[12]/data_i[24] ) );
  AO22X1_RVT U4111 ( .A1(\read_value_mux[12][25] ), .A2(n3025), .A3(
        write_data[25]), .A4(n3024), .Y(\words[12]/data_i[25] ) );
  AO22X1_RVT U4112 ( .A1(\read_value_mux[12][26] ), .A2(n3025), .A3(
        write_data[26]), .A4(n3024), .Y(\words[12]/data_i[26] ) );
  AO22X1_RVT U4113 ( .A1(\read_value_mux[12][27] ), .A2(n3025), .A3(
        write_data[27]), .A4(n3024), .Y(\words[12]/data_i[27] ) );
  AO22X1_RVT U4114 ( .A1(\read_value_mux[12][28] ), .A2(n3025), .A3(
        write_data[28]), .A4(n3024), .Y(\words[12]/data_i[28] ) );
  AO22X1_RVT U4115 ( .A1(\read_value_mux[12][29] ), .A2(n3025), .A3(
        write_data[29]), .A4(n3024), .Y(\words[12]/data_i[29] ) );
  AO22X1_RVT U4116 ( .A1(\read_value_mux[12][2] ), .A2(n3025), .A3(
        write_data[2]), .A4(n3024), .Y(\words[12]/data_i[2] ) );
  AO22X1_RVT U4117 ( .A1(n3024), .A2(write_data[30]), .A3(
        \read_value_mux[12][30] ), .A4(n3025), .Y(\words[12]/data_i[30] ) );
  AO22X1_RVT U4118 ( .A1(\read_value_mux[12][31] ), .A2(n3025), .A3(
        write_data[31]), .A4(n3024), .Y(\words[12]/data_i[31] ) );
  AO22X1_RVT U4119 ( .A1(\read_value_mux[12][3] ), .A2(n3025), .A3(
        write_data[3]), .A4(n3024), .Y(\words[12]/data_i[3] ) );
  AO22X1_RVT U4120 ( .A1(\read_value_mux[12][4] ), .A2(n3025), .A3(
        write_data[4]), .A4(n3024), .Y(\words[12]/data_i[4] ) );
  AO22X1_RVT U4121 ( .A1(\read_value_mux[12][5] ), .A2(n3025), .A3(
        write_data[5]), .A4(n3024), .Y(\words[12]/data_i[5] ) );
  AO22X1_RVT U4122 ( .A1(\read_value_mux[12][6] ), .A2(n3025), .A3(
        write_data[6]), .A4(n3024), .Y(\words[12]/data_i[6] ) );
  AO22X1_RVT U4123 ( .A1(\read_value_mux[12][7] ), .A2(n3025), .A3(
        write_data[7]), .A4(n3024), .Y(\words[12]/data_i[7] ) );
  AO22X1_RVT U4124 ( .A1(\read_value_mux[12][8] ), .A2(n3025), .A3(
        write_data[8]), .A4(n3024), .Y(\words[12]/data_i[8] ) );
  AO22X1_RVT U4125 ( .A1(\read_value_mux[12][9] ), .A2(n3025), .A3(
        write_data[9]), .A4(n3024), .Y(\words[12]/data_i[9] ) );
  AO21X1_RVT U4126 ( .A1(\words[12]/valid_o ), .A2(n3025), .A3(n3024), .Y(
        \words[12]/valid_i ) );
  AO22X1_RVT U4127 ( .A1(\read_value_mux[13][0] ), .A2(n1630), .A3(
        write_data[0]), .A4(n3028), .Y(\words[13]/data_i[0] ) );
  AO22X1_RVT U4128 ( .A1(\read_value_mux[13][10] ), .A2(n1630), .A3(
        write_data[10]), .A4(n3028), .Y(\words[13]/data_i[10] ) );
  AO22X1_RVT U4129 ( .A1(\read_value_mux[13][11] ), .A2(n1630), .A3(
        write_data[11]), .A4(n3028), .Y(\words[13]/data_i[11] ) );
  AO22X1_RVT U4130 ( .A1(\read_value_mux[13][12] ), .A2(n1630), .A3(
        write_data[12]), .A4(n3028), .Y(\words[13]/data_i[12] ) );
  AO22X1_RVT U4131 ( .A1(\read_value_mux[13][13] ), .A2(n1630), .A3(
        write_data[13]), .A4(n3028), .Y(\words[13]/data_i[13] ) );
  AO22X1_RVT U4132 ( .A1(\read_value_mux[13][14] ), .A2(n1630), .A3(
        write_data[14]), .A4(n3028), .Y(\words[13]/data_i[14] ) );
  AO22X1_RVT U4133 ( .A1(\read_value_mux[13][15] ), .A2(n1630), .A3(
        write_data[15]), .A4(n3028), .Y(\words[13]/data_i[15] ) );
  AO22X1_RVT U4134 ( .A1(\read_value_mux[13][16] ), .A2(n1630), .A3(
        write_data[16]), .A4(n3028), .Y(\words[13]/data_i[16] ) );
  AO22X1_RVT U4135 ( .A1(\read_value_mux[13][17] ), .A2(n1630), .A3(
        write_data[17]), .A4(n3028), .Y(\words[13]/data_i[17] ) );
  AO22X1_RVT U4136 ( .A1(\read_value_mux[13][18] ), .A2(n1630), .A3(
        write_data[18]), .A4(n3028), .Y(\words[13]/data_i[18] ) );
  AO22X1_RVT U4137 ( .A1(\read_value_mux[13][19] ), .A2(n1630), .A3(
        write_data[19]), .A4(n3028), .Y(\words[13]/data_i[19] ) );
  AO22X1_RVT U4138 ( .A1(n3028), .A2(write_data[1]), .A3(
        \read_value_mux[13][1] ), .A4(n1630), .Y(\words[13]/data_i[1] ) );
  AO22X1_RVT U4139 ( .A1(\read_value_mux[13][20] ), .A2(n1630), .A3(
        write_data[20]), .A4(n3028), .Y(\words[13]/data_i[20] ) );
  AO22X1_RVT U4140 ( .A1(\read_value_mux[13][21] ), .A2(n1630), .A3(
        write_data[21]), .A4(n3028), .Y(\words[13]/data_i[21] ) );
  AO22X1_RVT U4141 ( .A1(\read_value_mux[13][22] ), .A2(n1630), .A3(
        write_data[22]), .A4(n3028), .Y(\words[13]/data_i[22] ) );
  AO22X1_RVT U4142 ( .A1(\read_value_mux[13][23] ), .A2(n1630), .A3(
        write_data[23]), .A4(n3028), .Y(\words[13]/data_i[23] ) );
  AO22X1_RVT U4143 ( .A1(\read_value_mux[13][24] ), .A2(n1630), .A3(
        write_data[24]), .A4(n3028), .Y(\words[13]/data_i[24] ) );
  AO22X1_RVT U4144 ( .A1(\read_value_mux[13][25] ), .A2(n1630), .A3(
        write_data[25]), .A4(n3028), .Y(\words[13]/data_i[25] ) );
  AO22X1_RVT U4145 ( .A1(\read_value_mux[13][26] ), .A2(n1630), .A3(
        write_data[26]), .A4(n3028), .Y(\words[13]/data_i[26] ) );
  AO22X1_RVT U4146 ( .A1(\read_value_mux[13][27] ), .A2(n1630), .A3(
        write_data[27]), .A4(n3028), .Y(\words[13]/data_i[27] ) );
  AO22X1_RVT U4147 ( .A1(\read_value_mux[13][28] ), .A2(n1630), .A3(
        write_data[28]), .A4(n3028), .Y(\words[13]/data_i[28] ) );
  AO22X1_RVT U4148 ( .A1(\read_value_mux[13][29] ), .A2(n1630), .A3(
        write_data[29]), .A4(n3028), .Y(\words[13]/data_i[29] ) );
  AO22X1_RVT U4149 ( .A1(\read_value_mux[13][2] ), .A2(n1630), .A3(
        write_data[2]), .A4(n3028), .Y(\words[13]/data_i[2] ) );
  AO22X1_RVT U4150 ( .A1(n3028), .A2(write_data[30]), .A3(
        \read_value_mux[13][30] ), .A4(n1630), .Y(\words[13]/data_i[30] ) );
  AO22X1_RVT U4151 ( .A1(\read_value_mux[13][31] ), .A2(n1630), .A3(
        write_data[31]), .A4(n3028), .Y(\words[13]/data_i[31] ) );
  AO22X1_RVT U4152 ( .A1(\read_value_mux[13][3] ), .A2(n1630), .A3(
        write_data[3]), .A4(n3028), .Y(\words[13]/data_i[3] ) );
  AO22X1_RVT U4153 ( .A1(\read_value_mux[13][4] ), .A2(n1630), .A3(
        write_data[4]), .A4(n3028), .Y(\words[13]/data_i[4] ) );
  AO22X1_RVT U4154 ( .A1(\read_value_mux[13][5] ), .A2(n1630), .A3(
        write_data[5]), .A4(n3028), .Y(\words[13]/data_i[5] ) );
  AO22X1_RVT U4155 ( .A1(\read_value_mux[13][6] ), .A2(n1630), .A3(
        write_data[6]), .A4(n3028), .Y(\words[13]/data_i[6] ) );
  AO22X1_RVT U4156 ( .A1(\read_value_mux[13][7] ), .A2(n1630), .A3(
        write_data[7]), .A4(n3028), .Y(\words[13]/data_i[7] ) );
  AO22X1_RVT U4157 ( .A1(\read_value_mux[13][8] ), .A2(n1630), .A3(
        write_data[8]), .A4(n3028), .Y(\words[13]/data_i[8] ) );
  AO22X1_RVT U4158 ( .A1(\read_value_mux[13][9] ), .A2(n1630), .A3(
        write_data[9]), .A4(n3028), .Y(\words[13]/data_i[9] ) );
  AO21X1_RVT U4159 ( .A1(\words[13]/valid_o ), .A2(n1630), .A3(n3028), .Y(
        \words[13]/valid_i ) );
  AO22X1_RVT U4160 ( .A1(\read_value_mux[14][0] ), .A2(n3030), .A3(
        write_data[0]), .A4(n3029), .Y(\words[14]/data_i[0] ) );
  AO22X1_RVT U4161 ( .A1(\read_value_mux[14][10] ), .A2(n3030), .A3(
        write_data[10]), .A4(n3029), .Y(\words[14]/data_i[10] ) );
  AO22X1_RVT U4162 ( .A1(\read_value_mux[14][11] ), .A2(n3030), .A3(
        write_data[11]), .A4(n3029), .Y(\words[14]/data_i[11] ) );
  AO22X1_RVT U4163 ( .A1(\read_value_mux[14][12] ), .A2(n3030), .A3(
        write_data[12]), .A4(n3029), .Y(\words[14]/data_i[12] ) );
  AO22X1_RVT U4164 ( .A1(\read_value_mux[14][13] ), .A2(n3030), .A3(
        write_data[13]), .A4(n3029), .Y(\words[14]/data_i[13] ) );
  AO22X1_RVT U4165 ( .A1(\read_value_mux[14][14] ), .A2(n3030), .A3(
        write_data[14]), .A4(n3029), .Y(\words[14]/data_i[14] ) );
  AO22X1_RVT U4166 ( .A1(\read_value_mux[14][15] ), .A2(n3030), .A3(
        write_data[15]), .A4(n3029), .Y(\words[14]/data_i[15] ) );
  AO22X1_RVT U4167 ( .A1(\read_value_mux[14][16] ), .A2(n3030), .A3(
        write_data[16]), .A4(n3029), .Y(\words[14]/data_i[16] ) );
  AO22X1_RVT U4168 ( .A1(\read_value_mux[14][17] ), .A2(n3030), .A3(
        write_data[17]), .A4(n3029), .Y(\words[14]/data_i[17] ) );
  AO22X1_RVT U4169 ( .A1(\read_value_mux[14][18] ), .A2(n3030), .A3(
        write_data[18]), .A4(n3029), .Y(\words[14]/data_i[18] ) );
  AO22X1_RVT U4170 ( .A1(\read_value_mux[14][19] ), .A2(n3030), .A3(
        write_data[19]), .A4(n3029), .Y(\words[14]/data_i[19] ) );
  AO22X1_RVT U4171 ( .A1(n3029), .A2(write_data[1]), .A3(
        \read_value_mux[14][1] ), .A4(n3030), .Y(\words[14]/data_i[1] ) );
  AO22X1_RVT U4172 ( .A1(\read_value_mux[14][20] ), .A2(n3030), .A3(
        write_data[20]), .A4(n3029), .Y(\words[14]/data_i[20] ) );
  AO22X1_RVT U4173 ( .A1(\read_value_mux[14][21] ), .A2(n3030), .A3(
        write_data[21]), .A4(n3029), .Y(\words[14]/data_i[21] ) );
  AO22X1_RVT U4174 ( .A1(\read_value_mux[14][22] ), .A2(n3030), .A3(
        write_data[22]), .A4(n3029), .Y(\words[14]/data_i[22] ) );
  AO22X1_RVT U4175 ( .A1(\read_value_mux[14][23] ), .A2(n3030), .A3(
        write_data[23]), .A4(n3029), .Y(\words[14]/data_i[23] ) );
  AO22X1_RVT U4176 ( .A1(\read_value_mux[14][24] ), .A2(n3030), .A3(
        write_data[24]), .A4(n3029), .Y(\words[14]/data_i[24] ) );
  AO22X1_RVT U4177 ( .A1(\read_value_mux[14][25] ), .A2(n3030), .A3(
        write_data[25]), .A4(n3029), .Y(\words[14]/data_i[25] ) );
  AO22X1_RVT U4178 ( .A1(\read_value_mux[14][26] ), .A2(n3030), .A3(
        write_data[26]), .A4(n3029), .Y(\words[14]/data_i[26] ) );
  AO22X1_RVT U4179 ( .A1(\read_value_mux[14][27] ), .A2(n3030), .A3(
        write_data[27]), .A4(n3029), .Y(\words[14]/data_i[27] ) );
  AO22X1_RVT U4180 ( .A1(\read_value_mux[14][28] ), .A2(n3030), .A3(
        write_data[28]), .A4(n3029), .Y(\words[14]/data_i[28] ) );
  AO22X1_RVT U4181 ( .A1(\read_value_mux[14][29] ), .A2(n3030), .A3(
        write_data[29]), .A4(n3029), .Y(\words[14]/data_i[29] ) );
  AO22X1_RVT U4182 ( .A1(\read_value_mux[14][2] ), .A2(n3030), .A3(
        write_data[2]), .A4(n3029), .Y(\words[14]/data_i[2] ) );
  AO22X1_RVT U4183 ( .A1(n3029), .A2(write_data[30]), .A3(
        \read_value_mux[14][30] ), .A4(n3030), .Y(\words[14]/data_i[30] ) );
  AO22X1_RVT U4184 ( .A1(\read_value_mux[14][31] ), .A2(n3030), .A3(
        write_data[31]), .A4(n3029), .Y(\words[14]/data_i[31] ) );
  AO22X1_RVT U4185 ( .A1(\read_value_mux[14][3] ), .A2(n3030), .A3(
        write_data[3]), .A4(n3029), .Y(\words[14]/data_i[3] ) );
  AO22X1_RVT U4186 ( .A1(\read_value_mux[14][4] ), .A2(n3030), .A3(
        write_data[4]), .A4(n3029), .Y(\words[14]/data_i[4] ) );
  AO22X1_RVT U4187 ( .A1(\read_value_mux[14][5] ), .A2(n3030), .A3(
        write_data[5]), .A4(n3029), .Y(\words[14]/data_i[5] ) );
  AO22X1_RVT U4188 ( .A1(\read_value_mux[14][6] ), .A2(n3030), .A3(
        write_data[6]), .A4(n3029), .Y(\words[14]/data_i[6] ) );
  AO22X1_RVT U4189 ( .A1(\read_value_mux[14][7] ), .A2(n3030), .A3(
        write_data[7]), .A4(n3029), .Y(\words[14]/data_i[7] ) );
  AO22X1_RVT U4190 ( .A1(\read_value_mux[14][8] ), .A2(n3030), .A3(
        write_data[8]), .A4(n3029), .Y(\words[14]/data_i[8] ) );
  AO22X1_RVT U4191 ( .A1(\read_value_mux[14][9] ), .A2(n3030), .A3(
        write_data[9]), .A4(n3029), .Y(\words[14]/data_i[9] ) );
  AO21X1_RVT U4192 ( .A1(\words[14]/valid_o ), .A2(n3030), .A3(n3029), .Y(
        \words[14]/valid_i ) );
  AO22X1_RVT U4193 ( .A1(\read_value_mux[15][0] ), .A2(n1631), .A3(
        write_data[0]), .A4(n3033), .Y(\words[15]/data_i[0] ) );
  AO22X1_RVT U4194 ( .A1(\read_value_mux[15][10] ), .A2(n1631), .A3(
        write_data[10]), .A4(n3033), .Y(\words[15]/data_i[10] ) );
  AO22X1_RVT U4195 ( .A1(\read_value_mux[15][11] ), .A2(n1631), .A3(
        write_data[11]), .A4(n3033), .Y(\words[15]/data_i[11] ) );
  AO22X1_RVT U4196 ( .A1(\read_value_mux[15][12] ), .A2(n1631), .A3(
        write_data[12]), .A4(n3033), .Y(\words[15]/data_i[12] ) );
  AO22X1_RVT U4197 ( .A1(\read_value_mux[15][13] ), .A2(n1631), .A3(
        write_data[13]), .A4(n3033), .Y(\words[15]/data_i[13] ) );
  AO22X1_RVT U4198 ( .A1(\read_value_mux[15][14] ), .A2(n1631), .A3(
        write_data[14]), .A4(n3033), .Y(\words[15]/data_i[14] ) );
  AO22X1_RVT U4199 ( .A1(\read_value_mux[15][15] ), .A2(n1631), .A3(
        write_data[15]), .A4(n3033), .Y(\words[15]/data_i[15] ) );
  AO22X1_RVT U4200 ( .A1(\read_value_mux[15][16] ), .A2(n1631), .A3(
        write_data[16]), .A4(n3033), .Y(\words[15]/data_i[16] ) );
  AO22X1_RVT U4201 ( .A1(\read_value_mux[15][17] ), .A2(n1631), .A3(
        write_data[17]), .A4(n3033), .Y(\words[15]/data_i[17] ) );
  AO22X1_RVT U4202 ( .A1(\read_value_mux[15][18] ), .A2(n1631), .A3(
        write_data[18]), .A4(n3033), .Y(\words[15]/data_i[18] ) );
  AO22X1_RVT U4203 ( .A1(\read_value_mux[15][19] ), .A2(n1631), .A3(
        write_data[19]), .A4(n3033), .Y(\words[15]/data_i[19] ) );
  AO22X1_RVT U4204 ( .A1(n3033), .A2(write_data[1]), .A3(
        \read_value_mux[15][1] ), .A4(n1631), .Y(\words[15]/data_i[1] ) );
  AO22X1_RVT U4205 ( .A1(\read_value_mux[15][20] ), .A2(n1631), .A3(
        write_data[20]), .A4(n3033), .Y(\words[15]/data_i[20] ) );
  AO22X1_RVT U4206 ( .A1(\read_value_mux[15][21] ), .A2(n1631), .A3(
        write_data[21]), .A4(n3033), .Y(\words[15]/data_i[21] ) );
  AO22X1_RVT U4207 ( .A1(\read_value_mux[15][22] ), .A2(n1631), .A3(
        write_data[22]), .A4(n3033), .Y(\words[15]/data_i[22] ) );
  AO22X1_RVT U4208 ( .A1(\read_value_mux[15][23] ), .A2(n1631), .A3(
        write_data[23]), .A4(n3033), .Y(\words[15]/data_i[23] ) );
  AO22X1_RVT U4209 ( .A1(\read_value_mux[15][24] ), .A2(n1631), .A3(
        write_data[24]), .A4(n3033), .Y(\words[15]/data_i[24] ) );
  AO22X1_RVT U4210 ( .A1(\read_value_mux[15][25] ), .A2(n1631), .A3(
        write_data[25]), .A4(n3033), .Y(\words[15]/data_i[25] ) );
  AO22X1_RVT U4211 ( .A1(\read_value_mux[15][26] ), .A2(n1631), .A3(
        write_data[26]), .A4(n3033), .Y(\words[15]/data_i[26] ) );
  AO22X1_RVT U4212 ( .A1(\read_value_mux[15][27] ), .A2(n1631), .A3(
        write_data[27]), .A4(n3033), .Y(\words[15]/data_i[27] ) );
  AO22X1_RVT U4213 ( .A1(\read_value_mux[15][28] ), .A2(n1631), .A3(
        write_data[28]), .A4(n3033), .Y(\words[15]/data_i[28] ) );
  AO22X1_RVT U4214 ( .A1(\read_value_mux[15][29] ), .A2(n1631), .A3(
        write_data[29]), .A4(n3033), .Y(\words[15]/data_i[29] ) );
  AO22X1_RVT U4215 ( .A1(\read_value_mux[15][2] ), .A2(n1631), .A3(
        write_data[2]), .A4(n3033), .Y(\words[15]/data_i[2] ) );
  AO22X1_RVT U4216 ( .A1(n3033), .A2(write_data[30]), .A3(
        \read_value_mux[15][30] ), .A4(n1631), .Y(\words[15]/data_i[30] ) );
  AO22X1_RVT U4217 ( .A1(\read_value_mux[15][31] ), .A2(n1631), .A3(
        write_data[31]), .A4(n3033), .Y(\words[15]/data_i[31] ) );
  AO22X1_RVT U4218 ( .A1(\read_value_mux[15][3] ), .A2(n1631), .A3(
        write_data[3]), .A4(n3033), .Y(\words[15]/data_i[3] ) );
  AO22X1_RVT U4219 ( .A1(\read_value_mux[15][4] ), .A2(n1631), .A3(
        write_data[4]), .A4(n3033), .Y(\words[15]/data_i[4] ) );
  AO22X1_RVT U4220 ( .A1(\read_value_mux[15][5] ), .A2(n1631), .A3(
        write_data[5]), .A4(n3033), .Y(\words[15]/data_i[5] ) );
  AO22X1_RVT U4221 ( .A1(\read_value_mux[15][6] ), .A2(n1631), .A3(
        write_data[6]), .A4(n3033), .Y(\words[15]/data_i[6] ) );
  AO22X1_RVT U4222 ( .A1(\read_value_mux[15][7] ), .A2(n1631), .A3(
        write_data[7]), .A4(n3033), .Y(\words[15]/data_i[7] ) );
  AO22X1_RVT U4223 ( .A1(\read_value_mux[15][8] ), .A2(n1631), .A3(
        write_data[8]), .A4(n3033), .Y(\words[15]/data_i[8] ) );
  AO22X1_RVT U4224 ( .A1(\read_value_mux[15][9] ), .A2(n1631), .A3(
        write_data[9]), .A4(n3033), .Y(\words[15]/data_i[9] ) );
  AO21X1_RVT U4225 ( .A1(\words[15]/valid_o ), .A2(n1631), .A3(n3033), .Y(
        \words[15]/valid_i ) );
  NAND3X0_RVT U4226 ( .A1(write_index[4]), .A2(write), .A3(n3035), .Y(n3034)
         );
  AO22X1_RVT U4227 ( .A1(\read_value_mux[16][0] ), .A2(n1676), .A3(
        write_data[0]), .A4(n3036), .Y(\words[16]/data_i[0] ) );
  AO22X1_RVT U4228 ( .A1(\read_value_mux[16][10] ), .A2(n1676), .A3(
        write_data[10]), .A4(n3036), .Y(\words[16]/data_i[10] ) );
  AO22X1_RVT U4229 ( .A1(\read_value_mux[16][11] ), .A2(n1676), .A3(
        write_data[11]), .A4(n3036), .Y(\words[16]/data_i[11] ) );
  AO22X1_RVT U4230 ( .A1(\read_value_mux[16][12] ), .A2(n1676), .A3(
        write_data[12]), .A4(n3036), .Y(\words[16]/data_i[12] ) );
  AO22X1_RVT U4231 ( .A1(\read_value_mux[16][13] ), .A2(n1676), .A3(
        write_data[13]), .A4(n3036), .Y(\words[16]/data_i[13] ) );
  AO22X1_RVT U4232 ( .A1(\read_value_mux[16][14] ), .A2(n1676), .A3(
        write_data[14]), .A4(n3036), .Y(\words[16]/data_i[14] ) );
  AO22X1_RVT U4233 ( .A1(\read_value_mux[16][15] ), .A2(n1676), .A3(
        write_data[15]), .A4(n3036), .Y(\words[16]/data_i[15] ) );
  AO22X1_RVT U4234 ( .A1(\read_value_mux[16][16] ), .A2(n1676), .A3(
        write_data[16]), .A4(n3036), .Y(\words[16]/data_i[16] ) );
  AO22X1_RVT U4235 ( .A1(\read_value_mux[16][17] ), .A2(n1676), .A3(
        write_data[17]), .A4(n3036), .Y(\words[16]/data_i[17] ) );
  AO22X1_RVT U4236 ( .A1(\read_value_mux[16][18] ), .A2(n1676), .A3(
        write_data[18]), .A4(n3036), .Y(\words[16]/data_i[18] ) );
  AO22X1_RVT U4237 ( .A1(\read_value_mux[16][19] ), .A2(n1676), .A3(
        write_data[19]), .A4(n3036), .Y(\words[16]/data_i[19] ) );
  AO22X1_RVT U4238 ( .A1(n3036), .A2(write_data[1]), .A3(
        \read_value_mux[16][1] ), .A4(n1676), .Y(\words[16]/data_i[1] ) );
  AO22X1_RVT U4239 ( .A1(\read_value_mux[16][20] ), .A2(n1676), .A3(
        write_data[20]), .A4(n3036), .Y(\words[16]/data_i[20] ) );
  AO22X1_RVT U4240 ( .A1(\read_value_mux[16][21] ), .A2(n1676), .A3(
        write_data[21]), .A4(n3036), .Y(\words[16]/data_i[21] ) );
  AO22X1_RVT U4241 ( .A1(\read_value_mux[16][22] ), .A2(n1676), .A3(
        write_data[22]), .A4(n3036), .Y(\words[16]/data_i[22] ) );
  AO22X1_RVT U4242 ( .A1(\read_value_mux[16][23] ), .A2(n1676), .A3(
        write_data[23]), .A4(n3036), .Y(\words[16]/data_i[23] ) );
  AO22X1_RVT U4243 ( .A1(\read_value_mux[16][24] ), .A2(n1676), .A3(
        write_data[24]), .A4(n3036), .Y(\words[16]/data_i[24] ) );
  AO22X1_RVT U4244 ( .A1(\read_value_mux[16][25] ), .A2(n1676), .A3(
        write_data[25]), .A4(n3036), .Y(\words[16]/data_i[25] ) );
  AO22X1_RVT U4245 ( .A1(\read_value_mux[16][26] ), .A2(n1676), .A3(
        write_data[26]), .A4(n3036), .Y(\words[16]/data_i[26] ) );
  AO22X1_RVT U4246 ( .A1(\read_value_mux[16][27] ), .A2(n1676), .A3(
        write_data[27]), .A4(n3036), .Y(\words[16]/data_i[27] ) );
  AO22X1_RVT U4247 ( .A1(\read_value_mux[16][28] ), .A2(n1676), .A3(
        write_data[28]), .A4(n3036), .Y(\words[16]/data_i[28] ) );
  AO22X1_RVT U4248 ( .A1(\read_value_mux[16][29] ), .A2(n1676), .A3(
        write_data[29]), .A4(n3036), .Y(\words[16]/data_i[29] ) );
  AO22X1_RVT U4249 ( .A1(\read_value_mux[16][2] ), .A2(n1676), .A3(
        write_data[2]), .A4(n3036), .Y(\words[16]/data_i[2] ) );
  AO22X1_RVT U4250 ( .A1(n3036), .A2(write_data[30]), .A3(
        \read_value_mux[16][30] ), .A4(n1676), .Y(\words[16]/data_i[30] ) );
  AO22X1_RVT U4251 ( .A1(\read_value_mux[16][31] ), .A2(n1676), .A3(
        write_data[31]), .A4(n3036), .Y(\words[16]/data_i[31] ) );
  AO22X1_RVT U4252 ( .A1(\read_value_mux[16][3] ), .A2(n1676), .A3(
        write_data[3]), .A4(n3036), .Y(\words[16]/data_i[3] ) );
  AO22X1_RVT U4253 ( .A1(\read_value_mux[16][4] ), .A2(n1676), .A3(
        write_data[4]), .A4(n3036), .Y(\words[16]/data_i[4] ) );
  AO22X1_RVT U4254 ( .A1(\read_value_mux[16][5] ), .A2(n1676), .A3(
        write_data[5]), .A4(n3036), .Y(\words[16]/data_i[5] ) );
  AO22X1_RVT U4255 ( .A1(\read_value_mux[16][6] ), .A2(n1676), .A3(
        write_data[6]), .A4(n3036), .Y(\words[16]/data_i[6] ) );
  AO22X1_RVT U4256 ( .A1(\read_value_mux[16][7] ), .A2(n1676), .A3(
        write_data[7]), .A4(n3036), .Y(\words[16]/data_i[7] ) );
  AO22X1_RVT U4257 ( .A1(\read_value_mux[16][8] ), .A2(n1676), .A3(
        write_data[8]), .A4(n3036), .Y(\words[16]/data_i[8] ) );
  AO22X1_RVT U4258 ( .A1(\read_value_mux[16][9] ), .A2(n1676), .A3(
        write_data[9]), .A4(n3036), .Y(\words[16]/data_i[9] ) );
  AO21X1_RVT U4259 ( .A1(\words[16]/valid_o ), .A2(n1676), .A3(n3036), .Y(
        \words[16]/valid_i ) );
  AO22X1_RVT U4260 ( .A1(\read_value_mux[17][0] ), .A2(n1681), .A3(
        write_data[0]), .A4(n3037), .Y(\words[17]/data_i[0] ) );
  AO22X1_RVT U4261 ( .A1(\read_value_mux[17][10] ), .A2(n1681), .A3(
        write_data[10]), .A4(n3037), .Y(\words[17]/data_i[10] ) );
  AO22X1_RVT U4262 ( .A1(\read_value_mux[17][11] ), .A2(n1681), .A3(
        write_data[11]), .A4(n3037), .Y(\words[17]/data_i[11] ) );
  AO22X1_RVT U4263 ( .A1(\read_value_mux[17][12] ), .A2(n1681), .A3(
        write_data[12]), .A4(n3037), .Y(\words[17]/data_i[12] ) );
  AO22X1_RVT U4264 ( .A1(\read_value_mux[17][13] ), .A2(n1681), .A3(
        write_data[13]), .A4(n3037), .Y(\words[17]/data_i[13] ) );
  AO22X1_RVT U4265 ( .A1(\read_value_mux[17][14] ), .A2(n1681), .A3(
        write_data[14]), .A4(n3037), .Y(\words[17]/data_i[14] ) );
  AO22X1_RVT U4266 ( .A1(\read_value_mux[17][15] ), .A2(n1681), .A3(
        write_data[15]), .A4(n3037), .Y(\words[17]/data_i[15] ) );
  AO22X1_RVT U4267 ( .A1(\read_value_mux[17][16] ), .A2(n1681), .A3(
        write_data[16]), .A4(n3037), .Y(\words[17]/data_i[16] ) );
  AO22X1_RVT U4268 ( .A1(\read_value_mux[17][17] ), .A2(n1681), .A3(
        write_data[17]), .A4(n3037), .Y(\words[17]/data_i[17] ) );
  AO22X1_RVT U4269 ( .A1(\read_value_mux[17][18] ), .A2(n1681), .A3(
        write_data[18]), .A4(n3037), .Y(\words[17]/data_i[18] ) );
  AO22X1_RVT U4270 ( .A1(\read_value_mux[17][19] ), .A2(n1681), .A3(
        write_data[19]), .A4(n3037), .Y(\words[17]/data_i[19] ) );
  AO22X1_RVT U4271 ( .A1(n3037), .A2(write_data[1]), .A3(
        \read_value_mux[17][1] ), .A4(n1681), .Y(\words[17]/data_i[1] ) );
  AO22X1_RVT U4272 ( .A1(\read_value_mux[17][20] ), .A2(n1681), .A3(
        write_data[20]), .A4(n3037), .Y(\words[17]/data_i[20] ) );
  AO22X1_RVT U4273 ( .A1(\read_value_mux[17][21] ), .A2(n1681), .A3(
        write_data[21]), .A4(n3037), .Y(\words[17]/data_i[21] ) );
  AO22X1_RVT U4274 ( .A1(\read_value_mux[17][22] ), .A2(n1681), .A3(
        write_data[22]), .A4(n3037), .Y(\words[17]/data_i[22] ) );
  AO22X1_RVT U4275 ( .A1(\read_value_mux[17][23] ), .A2(n1681), .A3(
        write_data[23]), .A4(n3037), .Y(\words[17]/data_i[23] ) );
  AO22X1_RVT U4276 ( .A1(\read_value_mux[17][24] ), .A2(n1681), .A3(
        write_data[24]), .A4(n3037), .Y(\words[17]/data_i[24] ) );
  AO22X1_RVT U4277 ( .A1(\read_value_mux[17][25] ), .A2(n1681), .A3(
        write_data[25]), .A4(n3037), .Y(\words[17]/data_i[25] ) );
  AO22X1_RVT U4278 ( .A1(\read_value_mux[17][26] ), .A2(n1681), .A3(
        write_data[26]), .A4(n3037), .Y(\words[17]/data_i[26] ) );
  AO22X1_RVT U4279 ( .A1(\read_value_mux[17][27] ), .A2(n1681), .A3(
        write_data[27]), .A4(n3037), .Y(\words[17]/data_i[27] ) );
  AO22X1_RVT U4280 ( .A1(\read_value_mux[17][28] ), .A2(n1681), .A3(
        write_data[28]), .A4(n3037), .Y(\words[17]/data_i[28] ) );
  AO22X1_RVT U4281 ( .A1(\read_value_mux[17][29] ), .A2(n1681), .A3(
        write_data[29]), .A4(n3037), .Y(\words[17]/data_i[29] ) );
  AO22X1_RVT U4282 ( .A1(\read_value_mux[17][2] ), .A2(n1681), .A3(
        write_data[2]), .A4(n3037), .Y(\words[17]/data_i[2] ) );
  AO22X1_RVT U4283 ( .A1(n3037), .A2(write_data[30]), .A3(
        \read_value_mux[17][30] ), .A4(n1681), .Y(\words[17]/data_i[30] ) );
  AO22X1_RVT U4284 ( .A1(\read_value_mux[17][31] ), .A2(n1681), .A3(
        write_data[31]), .A4(n3037), .Y(\words[17]/data_i[31] ) );
  AO22X1_RVT U4285 ( .A1(\read_value_mux[17][3] ), .A2(n1681), .A3(
        write_data[3]), .A4(n3037), .Y(\words[17]/data_i[3] ) );
  AO22X1_RVT U4286 ( .A1(\read_value_mux[17][4] ), .A2(n1681), .A3(
        write_data[4]), .A4(n3037), .Y(\words[17]/data_i[4] ) );
  AO22X1_RVT U4287 ( .A1(\read_value_mux[17][5] ), .A2(n1681), .A3(
        write_data[5]), .A4(n3037), .Y(\words[17]/data_i[5] ) );
  AO22X1_RVT U4288 ( .A1(\read_value_mux[17][6] ), .A2(n1681), .A3(
        write_data[6]), .A4(n3037), .Y(\words[17]/data_i[6] ) );
  AO22X1_RVT U4289 ( .A1(\read_value_mux[17][7] ), .A2(n1681), .A3(
        write_data[7]), .A4(n3037), .Y(\words[17]/data_i[7] ) );
  AO22X1_RVT U4290 ( .A1(\read_value_mux[17][8] ), .A2(n1681), .A3(
        write_data[8]), .A4(n3037), .Y(\words[17]/data_i[8] ) );
  AO22X1_RVT U4291 ( .A1(\read_value_mux[17][9] ), .A2(n1681), .A3(
        write_data[9]), .A4(n3037), .Y(\words[17]/data_i[9] ) );
  AO21X1_RVT U4292 ( .A1(\words[17]/valid_o ), .A2(n1681), .A3(n3037), .Y(
        \words[17]/valid_i ) );
  AO22X1_RVT U4293 ( .A1(\read_value_mux[18][0] ), .A2(n3039), .A3(
        write_data[0]), .A4(n3038), .Y(\words[18]/data_i[0] ) );
  AO22X1_RVT U4294 ( .A1(\read_value_mux[18][10] ), .A2(n3039), .A3(
        write_data[10]), .A4(n3038), .Y(\words[18]/data_i[10] ) );
  AO22X1_RVT U4295 ( .A1(\read_value_mux[18][11] ), .A2(n3039), .A3(
        write_data[11]), .A4(n3038), .Y(\words[18]/data_i[11] ) );
  AO22X1_RVT U4296 ( .A1(\read_value_mux[18][12] ), .A2(n3039), .A3(
        write_data[12]), .A4(n3038), .Y(\words[18]/data_i[12] ) );
  AO22X1_RVT U4297 ( .A1(\read_value_mux[18][13] ), .A2(n3039), .A3(
        write_data[13]), .A4(n3038), .Y(\words[18]/data_i[13] ) );
  AO22X1_RVT U4298 ( .A1(\read_value_mux[18][14] ), .A2(n3039), .A3(
        write_data[14]), .A4(n3038), .Y(\words[18]/data_i[14] ) );
  AO22X1_RVT U4299 ( .A1(\read_value_mux[18][15] ), .A2(n3039), .A3(
        write_data[15]), .A4(n3038), .Y(\words[18]/data_i[15] ) );
  AO22X1_RVT U4300 ( .A1(\read_value_mux[18][16] ), .A2(n3039), .A3(
        write_data[16]), .A4(n3038), .Y(\words[18]/data_i[16] ) );
  AO22X1_RVT U4301 ( .A1(\read_value_mux[18][17] ), .A2(n3039), .A3(
        write_data[17]), .A4(n3038), .Y(\words[18]/data_i[17] ) );
  AO22X1_RVT U4302 ( .A1(\read_value_mux[18][18] ), .A2(n3039), .A3(
        write_data[18]), .A4(n3038), .Y(\words[18]/data_i[18] ) );
  AO22X1_RVT U4303 ( .A1(\read_value_mux[18][19] ), .A2(n3039), .A3(
        write_data[19]), .A4(n3038), .Y(\words[18]/data_i[19] ) );
  AO22X1_RVT U4304 ( .A1(n3038), .A2(write_data[1]), .A3(
        \read_value_mux[18][1] ), .A4(n3039), .Y(\words[18]/data_i[1] ) );
  AO22X1_RVT U4305 ( .A1(\read_value_mux[18][20] ), .A2(n3039), .A3(
        write_data[20]), .A4(n3038), .Y(\words[18]/data_i[20] ) );
  AO22X1_RVT U4306 ( .A1(\read_value_mux[18][21] ), .A2(n3039), .A3(
        write_data[21]), .A4(n3038), .Y(\words[18]/data_i[21] ) );
  AO22X1_RVT U4307 ( .A1(\read_value_mux[18][22] ), .A2(n3039), .A3(
        write_data[22]), .A4(n3038), .Y(\words[18]/data_i[22] ) );
  AO22X1_RVT U4308 ( .A1(\read_value_mux[18][23] ), .A2(n3039), .A3(
        write_data[23]), .A4(n3038), .Y(\words[18]/data_i[23] ) );
  AO22X1_RVT U4309 ( .A1(\read_value_mux[18][24] ), .A2(n3039), .A3(
        write_data[24]), .A4(n3038), .Y(\words[18]/data_i[24] ) );
  AO22X1_RVT U4310 ( .A1(\read_value_mux[18][25] ), .A2(n3039), .A3(
        write_data[25]), .A4(n3038), .Y(\words[18]/data_i[25] ) );
  AO22X1_RVT U4311 ( .A1(\read_value_mux[18][26] ), .A2(n3039), .A3(
        write_data[26]), .A4(n3038), .Y(\words[18]/data_i[26] ) );
  AO22X1_RVT U4312 ( .A1(\read_value_mux[18][27] ), .A2(n3039), .A3(
        write_data[27]), .A4(n3038), .Y(\words[18]/data_i[27] ) );
  AO22X1_RVT U4313 ( .A1(\read_value_mux[18][28] ), .A2(n3039), .A3(
        write_data[28]), .A4(n3038), .Y(\words[18]/data_i[28] ) );
  AO22X1_RVT U4314 ( .A1(\read_value_mux[18][29] ), .A2(n3039), .A3(
        write_data[29]), .A4(n3038), .Y(\words[18]/data_i[29] ) );
  AO22X1_RVT U4315 ( .A1(\read_value_mux[18][2] ), .A2(n3039), .A3(
        write_data[2]), .A4(n3038), .Y(\words[18]/data_i[2] ) );
  AO22X1_RVT U4316 ( .A1(n3038), .A2(write_data[30]), .A3(
        \read_value_mux[18][30] ), .A4(n3039), .Y(\words[18]/data_i[30] ) );
  AO22X1_RVT U4317 ( .A1(\read_value_mux[18][31] ), .A2(n3039), .A3(
        write_data[31]), .A4(n3038), .Y(\words[18]/data_i[31] ) );
  AO22X1_RVT U4318 ( .A1(\read_value_mux[18][3] ), .A2(n3039), .A3(
        write_data[3]), .A4(n3038), .Y(\words[18]/data_i[3] ) );
  AO22X1_RVT U4319 ( .A1(\read_value_mux[18][4] ), .A2(n3039), .A3(
        write_data[4]), .A4(n3038), .Y(\words[18]/data_i[4] ) );
  AO22X1_RVT U4320 ( .A1(\read_value_mux[18][5] ), .A2(n3039), .A3(
        write_data[5]), .A4(n3038), .Y(\words[18]/data_i[5] ) );
  AO22X1_RVT U4321 ( .A1(\read_value_mux[18][6] ), .A2(n3039), .A3(
        write_data[6]), .A4(n3038), .Y(\words[18]/data_i[6] ) );
  AO22X1_RVT U4322 ( .A1(\read_value_mux[18][7] ), .A2(n3039), .A3(
        write_data[7]), .A4(n3038), .Y(\words[18]/data_i[7] ) );
  AO22X1_RVT U4323 ( .A1(\read_value_mux[18][8] ), .A2(n3039), .A3(
        write_data[8]), .A4(n3038), .Y(\words[18]/data_i[8] ) );
  AO22X1_RVT U4324 ( .A1(\read_value_mux[18][9] ), .A2(n3039), .A3(
        write_data[9]), .A4(n3038), .Y(\words[18]/data_i[9] ) );
  AO21X1_RVT U4325 ( .A1(\words[18]/valid_o ), .A2(n3039), .A3(n3038), .Y(
        \words[18]/valid_i ) );
  AO22X1_RVT U4326 ( .A1(\read_value_mux[19][0] ), .A2(n3043), .A3(
        write_data[0]), .A4(n3042), .Y(\words[19]/data_i[0] ) );
  AO22X1_RVT U4327 ( .A1(\read_value_mux[19][10] ), .A2(n3043), .A3(
        write_data[10]), .A4(n3042), .Y(\words[19]/data_i[10] ) );
  AO22X1_RVT U4328 ( .A1(\read_value_mux[19][11] ), .A2(n3043), .A3(
        write_data[11]), .A4(n3042), .Y(\words[19]/data_i[11] ) );
  AO22X1_RVT U4329 ( .A1(\read_value_mux[19][12] ), .A2(n3043), .A3(
        write_data[12]), .A4(n3042), .Y(\words[19]/data_i[12] ) );
  AO22X1_RVT U4330 ( .A1(\read_value_mux[19][13] ), .A2(n3043), .A3(
        write_data[13]), .A4(n3042), .Y(\words[19]/data_i[13] ) );
  AO22X1_RVT U4331 ( .A1(\read_value_mux[19][14] ), .A2(n3043), .A3(
        write_data[14]), .A4(n3042), .Y(\words[19]/data_i[14] ) );
  AO22X1_RVT U4332 ( .A1(\read_value_mux[19][15] ), .A2(n3043), .A3(
        write_data[15]), .A4(n3042), .Y(\words[19]/data_i[15] ) );
  AO22X1_RVT U4333 ( .A1(\read_value_mux[19][16] ), .A2(n3043), .A3(
        write_data[16]), .A4(n3042), .Y(\words[19]/data_i[16] ) );
  AO22X1_RVT U4334 ( .A1(\read_value_mux[19][17] ), .A2(n3043), .A3(
        write_data[17]), .A4(n3042), .Y(\words[19]/data_i[17] ) );
  AO22X1_RVT U4335 ( .A1(\read_value_mux[19][18] ), .A2(n3043), .A3(
        write_data[18]), .A4(n3042), .Y(\words[19]/data_i[18] ) );
  AO22X1_RVT U4336 ( .A1(\read_value_mux[19][19] ), .A2(n3043), .A3(
        write_data[19]), .A4(n3042), .Y(\words[19]/data_i[19] ) );
  AO22X1_RVT U4337 ( .A1(n3042), .A2(write_data[1]), .A3(
        \read_value_mux[19][1] ), .A4(n3043), .Y(\words[19]/data_i[1] ) );
  AO22X1_RVT U4338 ( .A1(\read_value_mux[19][20] ), .A2(n3043), .A3(
        write_data[20]), .A4(n3042), .Y(\words[19]/data_i[20] ) );
  AO22X1_RVT U4339 ( .A1(\read_value_mux[19][21] ), .A2(n3043), .A3(
        write_data[21]), .A4(n3042), .Y(\words[19]/data_i[21] ) );
  AO22X1_RVT U4340 ( .A1(\read_value_mux[19][22] ), .A2(n3043), .A3(
        write_data[22]), .A4(n3042), .Y(\words[19]/data_i[22] ) );
  AO22X1_RVT U4341 ( .A1(\read_value_mux[19][23] ), .A2(n3043), .A3(
        write_data[23]), .A4(n3042), .Y(\words[19]/data_i[23] ) );
  AO22X1_RVT U4342 ( .A1(\read_value_mux[19][24] ), .A2(n3043), .A3(
        write_data[24]), .A4(n3042), .Y(\words[19]/data_i[24] ) );
  AO22X1_RVT U4343 ( .A1(\read_value_mux[19][25] ), .A2(n3043), .A3(
        write_data[25]), .A4(n3042), .Y(\words[19]/data_i[25] ) );
  AO22X1_RVT U4344 ( .A1(\read_value_mux[19][26] ), .A2(n3043), .A3(
        write_data[26]), .A4(n3042), .Y(\words[19]/data_i[26] ) );
  AO22X1_RVT U4345 ( .A1(\read_value_mux[19][27] ), .A2(n3043), .A3(
        write_data[27]), .A4(n3042), .Y(\words[19]/data_i[27] ) );
  AO22X1_RVT U4346 ( .A1(\read_value_mux[19][28] ), .A2(n3043), .A3(
        write_data[28]), .A4(n3042), .Y(\words[19]/data_i[28] ) );
  AO22X1_RVT U4347 ( .A1(\read_value_mux[19][29] ), .A2(n3043), .A3(
        write_data[29]), .A4(n3042), .Y(\words[19]/data_i[29] ) );
  AO22X1_RVT U4348 ( .A1(\read_value_mux[19][2] ), .A2(n3043), .A3(
        write_data[2]), .A4(n3042), .Y(\words[19]/data_i[2] ) );
  AO22X1_RVT U4349 ( .A1(n3042), .A2(write_data[30]), .A3(
        \read_value_mux[19][30] ), .A4(n3043), .Y(\words[19]/data_i[30] ) );
  AO22X1_RVT U4350 ( .A1(\read_value_mux[19][31] ), .A2(n3043), .A3(
        write_data[31]), .A4(n3042), .Y(\words[19]/data_i[31] ) );
  AO22X1_RVT U4351 ( .A1(\read_value_mux[19][3] ), .A2(n3043), .A3(
        write_data[3]), .A4(n3042), .Y(\words[19]/data_i[3] ) );
  AO22X1_RVT U4352 ( .A1(\read_value_mux[19][4] ), .A2(n3043), .A3(
        write_data[4]), .A4(n3042), .Y(\words[19]/data_i[4] ) );
  AO22X1_RVT U4353 ( .A1(\read_value_mux[19][5] ), .A2(n3043), .A3(
        write_data[5]), .A4(n3042), .Y(\words[19]/data_i[5] ) );
  AO22X1_RVT U4354 ( .A1(\read_value_mux[19][6] ), .A2(n3043), .A3(
        write_data[6]), .A4(n3042), .Y(\words[19]/data_i[6] ) );
  AO22X1_RVT U4355 ( .A1(\read_value_mux[19][7] ), .A2(n3043), .A3(
        write_data[7]), .A4(n3042), .Y(\words[19]/data_i[7] ) );
  AO22X1_RVT U4356 ( .A1(\read_value_mux[19][8] ), .A2(n3043), .A3(
        write_data[8]), .A4(n3042), .Y(\words[19]/data_i[8] ) );
  AO22X1_RVT U4357 ( .A1(\read_value_mux[19][9] ), .A2(n3043), .A3(
        write_data[9]), .A4(n3042), .Y(\words[19]/data_i[9] ) );
  AO21X1_RVT U4358 ( .A1(\words[19]/valid_o ), .A2(n3043), .A3(n3042), .Y(
        \words[19]/valid_i ) );
  AO22X1_RVT U4359 ( .A1(\read_value_mux[1][0] ), .A2(n1632), .A3(
        write_data[0]), .A4(n3044), .Y(\words[1]/data_i[0] ) );
  AO22X1_RVT U4360 ( .A1(\read_value_mux[1][10] ), .A2(n1632), .A3(
        write_data[10]), .A4(n3044), .Y(\words[1]/data_i[10] ) );
  AO22X1_RVT U4361 ( .A1(\read_value_mux[1][11] ), .A2(n1632), .A3(
        write_data[11]), .A4(n3044), .Y(\words[1]/data_i[11] ) );
  AO22X1_RVT U4362 ( .A1(\read_value_mux[1][12] ), .A2(n1632), .A3(
        write_data[12]), .A4(n3044), .Y(\words[1]/data_i[12] ) );
  AO22X1_RVT U4363 ( .A1(\read_value_mux[1][13] ), .A2(n1632), .A3(
        write_data[13]), .A4(n3044), .Y(\words[1]/data_i[13] ) );
  AO22X1_RVT U4364 ( .A1(\read_value_mux[1][14] ), .A2(n1632), .A3(
        write_data[14]), .A4(n3044), .Y(\words[1]/data_i[14] ) );
  AO22X1_RVT U4365 ( .A1(\read_value_mux[1][15] ), .A2(n1632), .A3(
        write_data[15]), .A4(n3044), .Y(\words[1]/data_i[15] ) );
  AO22X1_RVT U4366 ( .A1(\read_value_mux[1][16] ), .A2(n1632), .A3(
        write_data[16]), .A4(n3044), .Y(\words[1]/data_i[16] ) );
  AO22X1_RVT U4367 ( .A1(\read_value_mux[1][17] ), .A2(n1632), .A3(
        write_data[17]), .A4(n3044), .Y(\words[1]/data_i[17] ) );
  AO22X1_RVT U4368 ( .A1(\read_value_mux[1][18] ), .A2(n1632), .A3(
        write_data[18]), .A4(n3044), .Y(\words[1]/data_i[18] ) );
  AO22X1_RVT U4369 ( .A1(\read_value_mux[1][19] ), .A2(n1632), .A3(
        write_data[19]), .A4(n3044), .Y(\words[1]/data_i[19] ) );
  AO22X1_RVT U4370 ( .A1(n3044), .A2(write_data[1]), .A3(
        \read_value_mux[1][1] ), .A4(n1632), .Y(\words[1]/data_i[1] ) );
  AO22X1_RVT U4371 ( .A1(\read_value_mux[1][20] ), .A2(n1632), .A3(
        write_data[20]), .A4(n3044), .Y(\words[1]/data_i[20] ) );
  AO22X1_RVT U4372 ( .A1(\read_value_mux[1][21] ), .A2(n1632), .A3(
        write_data[21]), .A4(n3044), .Y(\words[1]/data_i[21] ) );
  AO22X1_RVT U4373 ( .A1(\read_value_mux[1][22] ), .A2(n1632), .A3(
        write_data[22]), .A4(n3044), .Y(\words[1]/data_i[22] ) );
  AO22X1_RVT U4374 ( .A1(\read_value_mux[1][23] ), .A2(n1632), .A3(
        write_data[23]), .A4(n3044), .Y(\words[1]/data_i[23] ) );
  AO22X1_RVT U4375 ( .A1(\read_value_mux[1][24] ), .A2(n1632), .A3(
        write_data[24]), .A4(n3044), .Y(\words[1]/data_i[24] ) );
  AO22X1_RVT U4376 ( .A1(\read_value_mux[1][25] ), .A2(n1632), .A3(
        write_data[25]), .A4(n3044), .Y(\words[1]/data_i[25] ) );
  AO22X1_RVT U4377 ( .A1(\read_value_mux[1][26] ), .A2(n1632), .A3(
        write_data[26]), .A4(n3044), .Y(\words[1]/data_i[26] ) );
  AO22X1_RVT U4378 ( .A1(\read_value_mux[1][27] ), .A2(n1632), .A3(
        write_data[27]), .A4(n3044), .Y(\words[1]/data_i[27] ) );
  AO22X1_RVT U4379 ( .A1(\read_value_mux[1][28] ), .A2(n1632), .A3(
        write_data[28]), .A4(n3044), .Y(\words[1]/data_i[28] ) );
  AO22X1_RVT U4380 ( .A1(\read_value_mux[1][29] ), .A2(n1632), .A3(
        write_data[29]), .A4(n3044), .Y(\words[1]/data_i[29] ) );
  AO22X1_RVT U4381 ( .A1(\read_value_mux[1][2] ), .A2(n1632), .A3(
        write_data[2]), .A4(n3044), .Y(\words[1]/data_i[2] ) );
  AO22X1_RVT U4382 ( .A1(n3044), .A2(write_data[30]), .A3(
        \read_value_mux[1][30] ), .A4(n1632), .Y(\words[1]/data_i[30] ) );
  AO22X1_RVT U4383 ( .A1(\read_value_mux[1][31] ), .A2(n1632), .A3(
        write_data[31]), .A4(n3044), .Y(\words[1]/data_i[31] ) );
  AO22X1_RVT U4384 ( .A1(\read_value_mux[1][3] ), .A2(n1632), .A3(
        write_data[3]), .A4(n3044), .Y(\words[1]/data_i[3] ) );
  AO22X1_RVT U4385 ( .A1(\read_value_mux[1][4] ), .A2(n1632), .A3(
        write_data[4]), .A4(n3044), .Y(\words[1]/data_i[4] ) );
  AO22X1_RVT U4386 ( .A1(\read_value_mux[1][5] ), .A2(n1632), .A3(
        write_data[5]), .A4(n3044), .Y(\words[1]/data_i[5] ) );
  AO22X1_RVT U4387 ( .A1(\read_value_mux[1][6] ), .A2(n1632), .A3(
        write_data[6]), .A4(n3044), .Y(\words[1]/data_i[6] ) );
  AO22X1_RVT U4388 ( .A1(\read_value_mux[1][7] ), .A2(n1632), .A3(
        write_data[7]), .A4(n3044), .Y(\words[1]/data_i[7] ) );
  AO22X1_RVT U4389 ( .A1(\read_value_mux[1][8] ), .A2(n1632), .A3(
        write_data[8]), .A4(n3044), .Y(\words[1]/data_i[8] ) );
  AO22X1_RVT U4390 ( .A1(\read_value_mux[1][9] ), .A2(n1632), .A3(
        write_data[9]), .A4(n3044), .Y(\words[1]/data_i[9] ) );
  AO21X1_RVT U4391 ( .A1(\words[1]/valid_o ), .A2(n1632), .A3(n3044), .Y(
        \words[1]/valid_i ) );
  AO22X1_RVT U4392 ( .A1(\read_value_mux[20][0] ), .A2(n3047), .A3(
        write_data[0]), .A4(n3046), .Y(\words[20]/data_i[0] ) );
  AO22X1_RVT U4393 ( .A1(\read_value_mux[20][10] ), .A2(n3047), .A3(
        write_data[10]), .A4(n3046), .Y(\words[20]/data_i[10] ) );
  AO22X1_RVT U4394 ( .A1(\read_value_mux[20][11] ), .A2(n3047), .A3(
        write_data[11]), .A4(n3046), .Y(\words[20]/data_i[11] ) );
  AO22X1_RVT U4395 ( .A1(\read_value_mux[20][12] ), .A2(n3047), .A3(
        write_data[12]), .A4(n3046), .Y(\words[20]/data_i[12] ) );
  AO22X1_RVT U4396 ( .A1(\read_value_mux[20][13] ), .A2(n3047), .A3(
        write_data[13]), .A4(n3046), .Y(\words[20]/data_i[13] ) );
  AO22X1_RVT U4397 ( .A1(\read_value_mux[20][14] ), .A2(n3047), .A3(
        write_data[14]), .A4(n3046), .Y(\words[20]/data_i[14] ) );
  AO22X1_RVT U4398 ( .A1(\read_value_mux[20][15] ), .A2(n3047), .A3(
        write_data[15]), .A4(n3046), .Y(\words[20]/data_i[15] ) );
  AO22X1_RVT U4399 ( .A1(\read_value_mux[20][16] ), .A2(n3047), .A3(
        write_data[16]), .A4(n3046), .Y(\words[20]/data_i[16] ) );
  AO22X1_RVT U4400 ( .A1(\read_value_mux[20][17] ), .A2(n3047), .A3(
        write_data[17]), .A4(n3046), .Y(\words[20]/data_i[17] ) );
  AO22X1_RVT U4401 ( .A1(\read_value_mux[20][18] ), .A2(n3047), .A3(
        write_data[18]), .A4(n3046), .Y(\words[20]/data_i[18] ) );
  AO22X1_RVT U4402 ( .A1(\read_value_mux[20][19] ), .A2(n3047), .A3(
        write_data[19]), .A4(n3046), .Y(\words[20]/data_i[19] ) );
  AO22X1_RVT U4403 ( .A1(n3046), .A2(write_data[1]), .A3(
        \read_value_mux[20][1] ), .A4(n3047), .Y(\words[20]/data_i[1] ) );
  AO22X1_RVT U4404 ( .A1(\read_value_mux[20][20] ), .A2(n3047), .A3(
        write_data[20]), .A4(n3046), .Y(\words[20]/data_i[20] ) );
  AO22X1_RVT U4405 ( .A1(\read_value_mux[20][21] ), .A2(n3047), .A3(
        write_data[21]), .A4(n3046), .Y(\words[20]/data_i[21] ) );
  AO22X1_RVT U4406 ( .A1(\read_value_mux[20][22] ), .A2(n3047), .A3(
        write_data[22]), .A4(n3046), .Y(\words[20]/data_i[22] ) );
  AO22X1_RVT U4407 ( .A1(\read_value_mux[20][23] ), .A2(n3047), .A3(
        write_data[23]), .A4(n3046), .Y(\words[20]/data_i[23] ) );
  AO22X1_RVT U4408 ( .A1(\read_value_mux[20][24] ), .A2(n3047), .A3(
        write_data[24]), .A4(n3046), .Y(\words[20]/data_i[24] ) );
  AO22X1_RVT U4409 ( .A1(\read_value_mux[20][25] ), .A2(n3047), .A3(
        write_data[25]), .A4(n3046), .Y(\words[20]/data_i[25] ) );
  AO22X1_RVT U4410 ( .A1(\read_value_mux[20][26] ), .A2(n3047), .A3(
        write_data[26]), .A4(n3046), .Y(\words[20]/data_i[26] ) );
  AO22X1_RVT U4411 ( .A1(\read_value_mux[20][27] ), .A2(n3047), .A3(
        write_data[27]), .A4(n3046), .Y(\words[20]/data_i[27] ) );
  AO22X1_RVT U4412 ( .A1(\read_value_mux[20][28] ), .A2(n3047), .A3(
        write_data[28]), .A4(n3046), .Y(\words[20]/data_i[28] ) );
  AO22X1_RVT U4413 ( .A1(\read_value_mux[20][29] ), .A2(n3047), .A3(
        write_data[29]), .A4(n3046), .Y(\words[20]/data_i[29] ) );
  AO22X1_RVT U4414 ( .A1(\read_value_mux[20][2] ), .A2(n3047), .A3(
        write_data[2]), .A4(n3046), .Y(\words[20]/data_i[2] ) );
  AO22X1_RVT U4415 ( .A1(n3046), .A2(write_data[30]), .A3(
        \read_value_mux[20][30] ), .A4(n3047), .Y(\words[20]/data_i[30] ) );
  AO22X1_RVT U4416 ( .A1(\read_value_mux[20][31] ), .A2(n3047), .A3(
        write_data[31]), .A4(n3046), .Y(\words[20]/data_i[31] ) );
  AO22X1_RVT U4417 ( .A1(\read_value_mux[20][3] ), .A2(n3047), .A3(
        write_data[3]), .A4(n3046), .Y(\words[20]/data_i[3] ) );
  AO22X1_RVT U4418 ( .A1(\read_value_mux[20][4] ), .A2(n3047), .A3(
        write_data[4]), .A4(n3046), .Y(\words[20]/data_i[4] ) );
  AO22X1_RVT U4419 ( .A1(\read_value_mux[20][5] ), .A2(n3047), .A3(
        write_data[5]), .A4(n3046), .Y(\words[20]/data_i[5] ) );
  AO22X1_RVT U4420 ( .A1(\read_value_mux[20][6] ), .A2(n3047), .A3(
        write_data[6]), .A4(n3046), .Y(\words[20]/data_i[6] ) );
  AO22X1_RVT U4421 ( .A1(\read_value_mux[20][7] ), .A2(n3047), .A3(
        write_data[7]), .A4(n3046), .Y(\words[20]/data_i[7] ) );
  AO22X1_RVT U4422 ( .A1(\read_value_mux[20][8] ), .A2(n3047), .A3(
        write_data[8]), .A4(n3046), .Y(\words[20]/data_i[8] ) );
  AO22X1_RVT U4423 ( .A1(\read_value_mux[20][9] ), .A2(n3047), .A3(
        write_data[9]), .A4(n3046), .Y(\words[20]/data_i[9] ) );
  AO21X1_RVT U4424 ( .A1(\words[20]/valid_o ), .A2(n3047), .A3(n3046), .Y(
        \words[20]/valid_i ) );
  AO22X1_RVT U4425 ( .A1(\read_value_mux[21][0] ), .A2(n1682), .A3(
        write_data[0]), .A4(n3048), .Y(\words[21]/data_i[0] ) );
  AO22X1_RVT U4426 ( .A1(\read_value_mux[21][10] ), .A2(n1682), .A3(
        write_data[10]), .A4(n3048), .Y(\words[21]/data_i[10] ) );
  AO22X1_RVT U4427 ( .A1(\read_value_mux[21][11] ), .A2(n1682), .A3(
        write_data[11]), .A4(n3048), .Y(\words[21]/data_i[11] ) );
  AO22X1_RVT U4428 ( .A1(\read_value_mux[21][12] ), .A2(n1682), .A3(
        write_data[12]), .A4(n3048), .Y(\words[21]/data_i[12] ) );
  AO22X1_RVT U4429 ( .A1(\read_value_mux[21][13] ), .A2(n1682), .A3(
        write_data[13]), .A4(n3048), .Y(\words[21]/data_i[13] ) );
  AO22X1_RVT U4430 ( .A1(\read_value_mux[21][14] ), .A2(n1682), .A3(
        write_data[14]), .A4(n3048), .Y(\words[21]/data_i[14] ) );
  AO22X1_RVT U4431 ( .A1(\read_value_mux[21][15] ), .A2(n1682), .A3(
        write_data[15]), .A4(n3048), .Y(\words[21]/data_i[15] ) );
  AO22X1_RVT U4432 ( .A1(\read_value_mux[21][16] ), .A2(n1682), .A3(
        write_data[16]), .A4(n3048), .Y(\words[21]/data_i[16] ) );
  AO22X1_RVT U4433 ( .A1(\read_value_mux[21][17] ), .A2(n1682), .A3(
        write_data[17]), .A4(n3048), .Y(\words[21]/data_i[17] ) );
  AO22X1_RVT U4434 ( .A1(\read_value_mux[21][18] ), .A2(n1682), .A3(
        write_data[18]), .A4(n3048), .Y(\words[21]/data_i[18] ) );
  AO22X1_RVT U4435 ( .A1(\read_value_mux[21][19] ), .A2(n1682), .A3(
        write_data[19]), .A4(n3048), .Y(\words[21]/data_i[19] ) );
  AO22X1_RVT U4436 ( .A1(n3048), .A2(write_data[1]), .A3(
        \read_value_mux[21][1] ), .A4(n1682), .Y(\words[21]/data_i[1] ) );
  AO22X1_RVT U4437 ( .A1(\read_value_mux[21][20] ), .A2(n1682), .A3(
        write_data[20]), .A4(n3048), .Y(\words[21]/data_i[20] ) );
  AO22X1_RVT U4438 ( .A1(\read_value_mux[21][21] ), .A2(n1682), .A3(
        write_data[21]), .A4(n3048), .Y(\words[21]/data_i[21] ) );
  AO22X1_RVT U4439 ( .A1(\read_value_mux[21][22] ), .A2(n1682), .A3(
        write_data[22]), .A4(n3048), .Y(\words[21]/data_i[22] ) );
  AO22X1_RVT U4440 ( .A1(\read_value_mux[21][23] ), .A2(n1682), .A3(
        write_data[23]), .A4(n3048), .Y(\words[21]/data_i[23] ) );
  AO22X1_RVT U4441 ( .A1(\read_value_mux[21][24] ), .A2(n1682), .A3(
        write_data[24]), .A4(n3048), .Y(\words[21]/data_i[24] ) );
  AO22X1_RVT U4442 ( .A1(\read_value_mux[21][25] ), .A2(n1682), .A3(
        write_data[25]), .A4(n3048), .Y(\words[21]/data_i[25] ) );
  AO22X1_RVT U4443 ( .A1(\read_value_mux[21][26] ), .A2(n1682), .A3(
        write_data[26]), .A4(n3048), .Y(\words[21]/data_i[26] ) );
  AO22X1_RVT U4444 ( .A1(\read_value_mux[21][27] ), .A2(n1682), .A3(
        write_data[27]), .A4(n3048), .Y(\words[21]/data_i[27] ) );
  AO22X1_RVT U4445 ( .A1(\read_value_mux[21][28] ), .A2(n1682), .A3(
        write_data[28]), .A4(n3048), .Y(\words[21]/data_i[28] ) );
  AO22X1_RVT U4446 ( .A1(\read_value_mux[21][29] ), .A2(n1682), .A3(
        write_data[29]), .A4(n3048), .Y(\words[21]/data_i[29] ) );
  AO22X1_RVT U4447 ( .A1(\read_value_mux[21][2] ), .A2(n1682), .A3(
        write_data[2]), .A4(n3048), .Y(\words[21]/data_i[2] ) );
  AO22X1_RVT U4448 ( .A1(n3048), .A2(write_data[30]), .A3(
        \read_value_mux[21][30] ), .A4(n1682), .Y(\words[21]/data_i[30] ) );
  AO22X1_RVT U4449 ( .A1(\read_value_mux[21][31] ), .A2(n1682), .A3(
        write_data[31]), .A4(n3048), .Y(\words[21]/data_i[31] ) );
  AO22X1_RVT U4450 ( .A1(\read_value_mux[21][3] ), .A2(n1682), .A3(
        write_data[3]), .A4(n3048), .Y(\words[21]/data_i[3] ) );
  AO22X1_RVT U4451 ( .A1(\read_value_mux[21][4] ), .A2(n1682), .A3(
        write_data[4]), .A4(n3048), .Y(\words[21]/data_i[4] ) );
  AO22X1_RVT U4452 ( .A1(\read_value_mux[21][5] ), .A2(n1682), .A3(
        write_data[5]), .A4(n3048), .Y(\words[21]/data_i[5] ) );
  AO22X1_RVT U4453 ( .A1(\read_value_mux[21][6] ), .A2(n1682), .A3(
        write_data[6]), .A4(n3048), .Y(\words[21]/data_i[6] ) );
  AO22X1_RVT U4454 ( .A1(\read_value_mux[21][7] ), .A2(n1682), .A3(
        write_data[7]), .A4(n3048), .Y(\words[21]/data_i[7] ) );
  AO22X1_RVT U4455 ( .A1(\read_value_mux[21][8] ), .A2(n1682), .A3(
        write_data[8]), .A4(n3048), .Y(\words[21]/data_i[8] ) );
  AO22X1_RVT U4456 ( .A1(\read_value_mux[21][9] ), .A2(n1682), .A3(
        write_data[9]), .A4(n3048), .Y(\words[21]/data_i[9] ) );
  AO21X1_RVT U4457 ( .A1(\words[21]/valid_o ), .A2(n1682), .A3(n3048), .Y(
        \words[21]/valid_i ) );
  AO22X1_RVT U4458 ( .A1(\read_value_mux[22][0] ), .A2(n3050), .A3(
        write_data[0]), .A4(n3049), .Y(\words[22]/data_i[0] ) );
  AO22X1_RVT U4459 ( .A1(\read_value_mux[22][10] ), .A2(n3050), .A3(
        write_data[10]), .A4(n3049), .Y(\words[22]/data_i[10] ) );
  AO22X1_RVT U4460 ( .A1(\read_value_mux[22][11] ), .A2(n3050), .A3(
        write_data[11]), .A4(n3049), .Y(\words[22]/data_i[11] ) );
  AO22X1_RVT U4461 ( .A1(\read_value_mux[22][12] ), .A2(n3050), .A3(
        write_data[12]), .A4(n3049), .Y(\words[22]/data_i[12] ) );
  AO22X1_RVT U4462 ( .A1(\read_value_mux[22][13] ), .A2(n3050), .A3(
        write_data[13]), .A4(n3049), .Y(\words[22]/data_i[13] ) );
  AO22X1_RVT U4463 ( .A1(\read_value_mux[22][14] ), .A2(n3050), .A3(
        write_data[14]), .A4(n3049), .Y(\words[22]/data_i[14] ) );
  AO22X1_RVT U4464 ( .A1(\read_value_mux[22][15] ), .A2(n3050), .A3(
        write_data[15]), .A4(n3049), .Y(\words[22]/data_i[15] ) );
  AO22X1_RVT U4465 ( .A1(\read_value_mux[22][16] ), .A2(n3050), .A3(
        write_data[16]), .A4(n3049), .Y(\words[22]/data_i[16] ) );
  AO22X1_RVT U4466 ( .A1(\read_value_mux[22][17] ), .A2(n3050), .A3(
        write_data[17]), .A4(n3049), .Y(\words[22]/data_i[17] ) );
  AO22X1_RVT U4467 ( .A1(\read_value_mux[22][18] ), .A2(n3050), .A3(
        write_data[18]), .A4(n3049), .Y(\words[22]/data_i[18] ) );
  AO22X1_RVT U4468 ( .A1(\read_value_mux[22][19] ), .A2(n3050), .A3(
        write_data[19]), .A4(n3049), .Y(\words[22]/data_i[19] ) );
  AO22X1_RVT U4469 ( .A1(n3049), .A2(write_data[1]), .A3(
        \read_value_mux[22][1] ), .A4(n3050), .Y(\words[22]/data_i[1] ) );
  AO22X1_RVT U4470 ( .A1(\read_value_mux[22][20] ), .A2(n3050), .A3(
        write_data[20]), .A4(n3049), .Y(\words[22]/data_i[20] ) );
  AO22X1_RVT U4471 ( .A1(\read_value_mux[22][21] ), .A2(n3050), .A3(
        write_data[21]), .A4(n3049), .Y(\words[22]/data_i[21] ) );
  AO22X1_RVT U4472 ( .A1(\read_value_mux[22][22] ), .A2(n3050), .A3(
        write_data[22]), .A4(n3049), .Y(\words[22]/data_i[22] ) );
  AO22X1_RVT U4473 ( .A1(\read_value_mux[22][23] ), .A2(n3050), .A3(
        write_data[23]), .A4(n3049), .Y(\words[22]/data_i[23] ) );
  AO22X1_RVT U4474 ( .A1(\read_value_mux[22][24] ), .A2(n3050), .A3(
        write_data[24]), .A4(n3049), .Y(\words[22]/data_i[24] ) );
  AO22X1_RVT U4475 ( .A1(\read_value_mux[22][25] ), .A2(n3050), .A3(
        write_data[25]), .A4(n3049), .Y(\words[22]/data_i[25] ) );
  AO22X1_RVT U4476 ( .A1(\read_value_mux[22][26] ), .A2(n3050), .A3(
        write_data[26]), .A4(n3049), .Y(\words[22]/data_i[26] ) );
  AO22X1_RVT U4477 ( .A1(\read_value_mux[22][27] ), .A2(n3050), .A3(
        write_data[27]), .A4(n3049), .Y(\words[22]/data_i[27] ) );
  AO22X1_RVT U4478 ( .A1(\read_value_mux[22][28] ), .A2(n3050), .A3(
        write_data[28]), .A4(n3049), .Y(\words[22]/data_i[28] ) );
  AO22X1_RVT U4479 ( .A1(\read_value_mux[22][29] ), .A2(n3050), .A3(
        write_data[29]), .A4(n3049), .Y(\words[22]/data_i[29] ) );
  AO22X1_RVT U4480 ( .A1(\read_value_mux[22][2] ), .A2(n3050), .A3(
        write_data[2]), .A4(n3049), .Y(\words[22]/data_i[2] ) );
  AO22X1_RVT U4481 ( .A1(n3049), .A2(write_data[30]), .A3(
        \read_value_mux[22][30] ), .A4(n3050), .Y(\words[22]/data_i[30] ) );
  AO22X1_RVT U4482 ( .A1(\read_value_mux[22][31] ), .A2(n3050), .A3(
        write_data[31]), .A4(n3049), .Y(\words[22]/data_i[31] ) );
  AO22X1_RVT U4483 ( .A1(\read_value_mux[22][3] ), .A2(n3050), .A3(
        write_data[3]), .A4(n3049), .Y(\words[22]/data_i[3] ) );
  AO22X1_RVT U4484 ( .A1(\read_value_mux[22][4] ), .A2(n3050), .A3(
        write_data[4]), .A4(n3049), .Y(\words[22]/data_i[4] ) );
  AO22X1_RVT U4485 ( .A1(\read_value_mux[22][5] ), .A2(n3050), .A3(
        write_data[5]), .A4(n3049), .Y(\words[22]/data_i[5] ) );
  AO22X1_RVT U4486 ( .A1(\read_value_mux[22][6] ), .A2(n3050), .A3(
        write_data[6]), .A4(n3049), .Y(\words[22]/data_i[6] ) );
  AO22X1_RVT U4487 ( .A1(\read_value_mux[22][7] ), .A2(n3050), .A3(
        write_data[7]), .A4(n3049), .Y(\words[22]/data_i[7] ) );
  AO22X1_RVT U4488 ( .A1(\read_value_mux[22][8] ), .A2(n3050), .A3(
        write_data[8]), .A4(n3049), .Y(\words[22]/data_i[8] ) );
  AO22X1_RVT U4489 ( .A1(\read_value_mux[22][9] ), .A2(n3050), .A3(
        write_data[9]), .A4(n3049), .Y(\words[22]/data_i[9] ) );
  AO21X1_RVT U4490 ( .A1(\words[22]/valid_o ), .A2(n3050), .A3(n3049), .Y(
        \words[22]/valid_i ) );
  AO22X1_RVT U4491 ( .A1(\read_value_mux[23][0] ), .A2(n3054), .A3(
        write_data[0]), .A4(n3053), .Y(\words[23]/data_i[0] ) );
  AO22X1_RVT U4492 ( .A1(\read_value_mux[23][10] ), .A2(n3054), .A3(
        write_data[10]), .A4(n3053), .Y(\words[23]/data_i[10] ) );
  AO22X1_RVT U4493 ( .A1(\read_value_mux[23][11] ), .A2(n3054), .A3(
        write_data[11]), .A4(n3053), .Y(\words[23]/data_i[11] ) );
  AO22X1_RVT U4494 ( .A1(\read_value_mux[23][12] ), .A2(n3054), .A3(
        write_data[12]), .A4(n3053), .Y(\words[23]/data_i[12] ) );
  AO22X1_RVT U4495 ( .A1(\read_value_mux[23][13] ), .A2(n3054), .A3(
        write_data[13]), .A4(n3053), .Y(\words[23]/data_i[13] ) );
  AO22X1_RVT U4496 ( .A1(\read_value_mux[23][14] ), .A2(n3054), .A3(
        write_data[14]), .A4(n3053), .Y(\words[23]/data_i[14] ) );
  AO22X1_RVT U4497 ( .A1(\read_value_mux[23][15] ), .A2(n3054), .A3(
        write_data[15]), .A4(n3053), .Y(\words[23]/data_i[15] ) );
  AO22X1_RVT U4498 ( .A1(\read_value_mux[23][16] ), .A2(n3054), .A3(
        write_data[16]), .A4(n3053), .Y(\words[23]/data_i[16] ) );
  AO22X1_RVT U4499 ( .A1(\read_value_mux[23][17] ), .A2(n3054), .A3(
        write_data[17]), .A4(n3053), .Y(\words[23]/data_i[17] ) );
  AO22X1_RVT U4500 ( .A1(\read_value_mux[23][18] ), .A2(n3054), .A3(
        write_data[18]), .A4(n3053), .Y(\words[23]/data_i[18] ) );
  AO22X1_RVT U4501 ( .A1(\read_value_mux[23][19] ), .A2(n3054), .A3(
        write_data[19]), .A4(n3053), .Y(\words[23]/data_i[19] ) );
  AO22X1_RVT U4502 ( .A1(n3053), .A2(write_data[1]), .A3(
        \read_value_mux[23][1] ), .A4(n3054), .Y(\words[23]/data_i[1] ) );
  AO22X1_RVT U4503 ( .A1(\read_value_mux[23][20] ), .A2(n3054), .A3(
        write_data[20]), .A4(n3053), .Y(\words[23]/data_i[20] ) );
  AO22X1_RVT U4504 ( .A1(\read_value_mux[23][21] ), .A2(n3054), .A3(
        write_data[21]), .A4(n3053), .Y(\words[23]/data_i[21] ) );
  AO22X1_RVT U4505 ( .A1(\read_value_mux[23][22] ), .A2(n3054), .A3(
        write_data[22]), .A4(n3053), .Y(\words[23]/data_i[22] ) );
  AO22X1_RVT U4506 ( .A1(\read_value_mux[23][23] ), .A2(n3054), .A3(
        write_data[23]), .A4(n3053), .Y(\words[23]/data_i[23] ) );
  AO22X1_RVT U4507 ( .A1(\read_value_mux[23][24] ), .A2(n3054), .A3(
        write_data[24]), .A4(n3053), .Y(\words[23]/data_i[24] ) );
  AO22X1_RVT U4508 ( .A1(\read_value_mux[23][25] ), .A2(n3054), .A3(
        write_data[25]), .A4(n3053), .Y(\words[23]/data_i[25] ) );
  AO22X1_RVT U4509 ( .A1(\read_value_mux[23][26] ), .A2(n3054), .A3(
        write_data[26]), .A4(n3053), .Y(\words[23]/data_i[26] ) );
  AO22X1_RVT U4510 ( .A1(\read_value_mux[23][27] ), .A2(n3054), .A3(
        write_data[27]), .A4(n3053), .Y(\words[23]/data_i[27] ) );
  AO22X1_RVT U4511 ( .A1(\read_value_mux[23][28] ), .A2(n3054), .A3(
        write_data[28]), .A4(n3053), .Y(\words[23]/data_i[28] ) );
  AO22X1_RVT U4512 ( .A1(\read_value_mux[23][29] ), .A2(n3054), .A3(
        write_data[29]), .A4(n3053), .Y(\words[23]/data_i[29] ) );
  AO22X1_RVT U4513 ( .A1(\read_value_mux[23][2] ), .A2(n3054), .A3(
        write_data[2]), .A4(n3053), .Y(\words[23]/data_i[2] ) );
  AO22X1_RVT U4514 ( .A1(n3053), .A2(write_data[30]), .A3(
        \read_value_mux[23][30] ), .A4(n3054), .Y(\words[23]/data_i[30] ) );
  AO22X1_RVT U4515 ( .A1(\read_value_mux[23][31] ), .A2(n3054), .A3(
        write_data[31]), .A4(n3053), .Y(\words[23]/data_i[31] ) );
  AO22X1_RVT U4516 ( .A1(\read_value_mux[23][3] ), .A2(n3054), .A3(
        write_data[3]), .A4(n3053), .Y(\words[23]/data_i[3] ) );
  AO22X1_RVT U4517 ( .A1(\read_value_mux[23][4] ), .A2(n3054), .A3(
        write_data[4]), .A4(n3053), .Y(\words[23]/data_i[4] ) );
  AO22X1_RVT U4518 ( .A1(\read_value_mux[23][5] ), .A2(n3054), .A3(
        write_data[5]), .A4(n3053), .Y(\words[23]/data_i[5] ) );
  AO22X1_RVT U4519 ( .A1(\read_value_mux[23][6] ), .A2(n3054), .A3(
        write_data[6]), .A4(n3053), .Y(\words[23]/data_i[6] ) );
  AO22X1_RVT U4520 ( .A1(\read_value_mux[23][7] ), .A2(n3054), .A3(
        write_data[7]), .A4(n3053), .Y(\words[23]/data_i[7] ) );
  AO22X1_RVT U4521 ( .A1(\read_value_mux[23][8] ), .A2(n3054), .A3(
        write_data[8]), .A4(n3053), .Y(\words[23]/data_i[8] ) );
  AO22X1_RVT U4522 ( .A1(\read_value_mux[23][9] ), .A2(n3054), .A3(
        write_data[9]), .A4(n3053), .Y(\words[23]/data_i[9] ) );
  AO21X1_RVT U4523 ( .A1(\words[23]/valid_o ), .A2(n3054), .A3(n3053), .Y(
        \words[23]/valid_i ) );
  AO22X1_RVT U4524 ( .A1(\read_value_mux[24][0] ), .A2(n1677), .A3(
        write_data[0]), .A4(n3055), .Y(\words[24]/data_i[0] ) );
  AO22X1_RVT U4525 ( .A1(\read_value_mux[24][10] ), .A2(n1677), .A3(
        write_data[10]), .A4(n3055), .Y(\words[24]/data_i[10] ) );
  AO22X1_RVT U4526 ( .A1(\read_value_mux[24][11] ), .A2(n1677), .A3(
        write_data[11]), .A4(n3055), .Y(\words[24]/data_i[11] ) );
  AO22X1_RVT U4527 ( .A1(\read_value_mux[24][12] ), .A2(n1677), .A3(
        write_data[12]), .A4(n3055), .Y(\words[24]/data_i[12] ) );
  AO22X1_RVT U4528 ( .A1(\read_value_mux[24][13] ), .A2(n1677), .A3(
        write_data[13]), .A4(n3055), .Y(\words[24]/data_i[13] ) );
  AO22X1_RVT U4529 ( .A1(\read_value_mux[24][14] ), .A2(n1677), .A3(
        write_data[14]), .A4(n3055), .Y(\words[24]/data_i[14] ) );
  AO22X1_RVT U4530 ( .A1(\read_value_mux[24][15] ), .A2(n1677), .A3(
        write_data[15]), .A4(n3055), .Y(\words[24]/data_i[15] ) );
  AO22X1_RVT U4531 ( .A1(\read_value_mux[24][16] ), .A2(n1677), .A3(
        write_data[16]), .A4(n3055), .Y(\words[24]/data_i[16] ) );
  AO22X1_RVT U4532 ( .A1(\read_value_mux[24][17] ), .A2(n1677), .A3(
        write_data[17]), .A4(n3055), .Y(\words[24]/data_i[17] ) );
  AO22X1_RVT U4533 ( .A1(\read_value_mux[24][18] ), .A2(n1677), .A3(
        write_data[18]), .A4(n3055), .Y(\words[24]/data_i[18] ) );
  AO22X1_RVT U4534 ( .A1(\read_value_mux[24][19] ), .A2(n1677), .A3(
        write_data[19]), .A4(n3055), .Y(\words[24]/data_i[19] ) );
  AO22X1_RVT U4535 ( .A1(n3055), .A2(write_data[1]), .A3(
        \read_value_mux[24][1] ), .A4(n1677), .Y(\words[24]/data_i[1] ) );
  AO22X1_RVT U4536 ( .A1(\read_value_mux[24][20] ), .A2(n1677), .A3(
        write_data[20]), .A4(n3055), .Y(\words[24]/data_i[20] ) );
  AO22X1_RVT U4537 ( .A1(\read_value_mux[24][21] ), .A2(n1677), .A3(
        write_data[21]), .A4(n3055), .Y(\words[24]/data_i[21] ) );
  AO22X1_RVT U4538 ( .A1(\read_value_mux[24][22] ), .A2(n1677), .A3(
        write_data[22]), .A4(n3055), .Y(\words[24]/data_i[22] ) );
  AO22X1_RVT U4539 ( .A1(\read_value_mux[24][23] ), .A2(n1677), .A3(
        write_data[23]), .A4(n3055), .Y(\words[24]/data_i[23] ) );
  AO22X1_RVT U4540 ( .A1(\read_value_mux[24][24] ), .A2(n1677), .A3(
        write_data[24]), .A4(n3055), .Y(\words[24]/data_i[24] ) );
  AO22X1_RVT U4541 ( .A1(\read_value_mux[24][25] ), .A2(n1677), .A3(
        write_data[25]), .A4(n3055), .Y(\words[24]/data_i[25] ) );
  AO22X1_RVT U4542 ( .A1(\read_value_mux[24][26] ), .A2(n1677), .A3(
        write_data[26]), .A4(n3055), .Y(\words[24]/data_i[26] ) );
  AO22X1_RVT U4543 ( .A1(\read_value_mux[24][27] ), .A2(n1677), .A3(
        write_data[27]), .A4(n3055), .Y(\words[24]/data_i[27] ) );
  AO22X1_RVT U4544 ( .A1(\read_value_mux[24][28] ), .A2(n1677), .A3(
        write_data[28]), .A4(n3055), .Y(\words[24]/data_i[28] ) );
  AO22X1_RVT U4545 ( .A1(\read_value_mux[24][29] ), .A2(n1677), .A3(
        write_data[29]), .A4(n3055), .Y(\words[24]/data_i[29] ) );
  AO22X1_RVT U4546 ( .A1(\read_value_mux[24][2] ), .A2(n1677), .A3(
        write_data[2]), .A4(n3055), .Y(\words[24]/data_i[2] ) );
  AO22X1_RVT U4547 ( .A1(n3055), .A2(write_data[30]), .A3(
        \read_value_mux[24][30] ), .A4(n1677), .Y(\words[24]/data_i[30] ) );
  AO22X1_RVT U4548 ( .A1(\read_value_mux[24][31] ), .A2(n1677), .A3(
        write_data[31]), .A4(n3055), .Y(\words[24]/data_i[31] ) );
  AO22X1_RVT U4549 ( .A1(\read_value_mux[24][3] ), .A2(n1677), .A3(
        write_data[3]), .A4(n3055), .Y(\words[24]/data_i[3] ) );
  AO22X1_RVT U4550 ( .A1(\read_value_mux[24][4] ), .A2(n1677), .A3(
        write_data[4]), .A4(n3055), .Y(\words[24]/data_i[4] ) );
  AO22X1_RVT U4551 ( .A1(\read_value_mux[24][5] ), .A2(n1677), .A3(
        write_data[5]), .A4(n3055), .Y(\words[24]/data_i[5] ) );
  AO22X1_RVT U4552 ( .A1(\read_value_mux[24][6] ), .A2(n1677), .A3(
        write_data[6]), .A4(n3055), .Y(\words[24]/data_i[6] ) );
  AO22X1_RVT U4553 ( .A1(\read_value_mux[24][7] ), .A2(n1677), .A3(
        write_data[7]), .A4(n3055), .Y(\words[24]/data_i[7] ) );
  AO22X1_RVT U4554 ( .A1(\read_value_mux[24][8] ), .A2(n1677), .A3(
        write_data[8]), .A4(n3055), .Y(\words[24]/data_i[8] ) );
  AO22X1_RVT U4555 ( .A1(\read_value_mux[24][9] ), .A2(n1677), .A3(
        write_data[9]), .A4(n3055), .Y(\words[24]/data_i[9] ) );
  AO21X1_RVT U4556 ( .A1(\words[24]/valid_o ), .A2(n1677), .A3(n3055), .Y(
        \words[24]/valid_i ) );
  AO22X1_RVT U4557 ( .A1(\read_value_mux[25][0] ), .A2(n1683), .A3(
        write_data[0]), .A4(n3056), .Y(\words[25]/data_i[0] ) );
  AO22X1_RVT U4558 ( .A1(\read_value_mux[25][10] ), .A2(n1683), .A3(
        write_data[10]), .A4(n3056), .Y(\words[25]/data_i[10] ) );
  AO22X1_RVT U4559 ( .A1(\read_value_mux[25][11] ), .A2(n1683), .A3(
        write_data[11]), .A4(n3056), .Y(\words[25]/data_i[11] ) );
  AO22X1_RVT U4560 ( .A1(\read_value_mux[25][12] ), .A2(n1683), .A3(
        write_data[12]), .A4(n3056), .Y(\words[25]/data_i[12] ) );
  AO22X1_RVT U4561 ( .A1(\read_value_mux[25][13] ), .A2(n1683), .A3(
        write_data[13]), .A4(n3056), .Y(\words[25]/data_i[13] ) );
  AO22X1_RVT U4562 ( .A1(\read_value_mux[25][14] ), .A2(n1683), .A3(
        write_data[14]), .A4(n3056), .Y(\words[25]/data_i[14] ) );
  AO22X1_RVT U4563 ( .A1(\read_value_mux[25][15] ), .A2(n1683), .A3(
        write_data[15]), .A4(n3056), .Y(\words[25]/data_i[15] ) );
  AO22X1_RVT U4564 ( .A1(\read_value_mux[25][16] ), .A2(n1683), .A3(
        write_data[16]), .A4(n3056), .Y(\words[25]/data_i[16] ) );
  AO22X1_RVT U4565 ( .A1(\read_value_mux[25][17] ), .A2(n1683), .A3(
        write_data[17]), .A4(n3056), .Y(\words[25]/data_i[17] ) );
  AO22X1_RVT U4566 ( .A1(\read_value_mux[25][18] ), .A2(n1683), .A3(
        write_data[18]), .A4(n3056), .Y(\words[25]/data_i[18] ) );
  AO22X1_RVT U4567 ( .A1(\read_value_mux[25][19] ), .A2(n1683), .A3(
        write_data[19]), .A4(n3056), .Y(\words[25]/data_i[19] ) );
  AO22X1_RVT U4568 ( .A1(n3056), .A2(write_data[1]), .A3(
        \read_value_mux[25][1] ), .A4(n1683), .Y(\words[25]/data_i[1] ) );
  AO22X1_RVT U4569 ( .A1(\read_value_mux[25][20] ), .A2(n1683), .A3(
        write_data[20]), .A4(n3056), .Y(\words[25]/data_i[20] ) );
  AO22X1_RVT U4570 ( .A1(\read_value_mux[25][21] ), .A2(n1683), .A3(
        write_data[21]), .A4(n3056), .Y(\words[25]/data_i[21] ) );
  AO22X1_RVT U4571 ( .A1(\read_value_mux[25][22] ), .A2(n1683), .A3(
        write_data[22]), .A4(n3056), .Y(\words[25]/data_i[22] ) );
  AO22X1_RVT U4572 ( .A1(\read_value_mux[25][23] ), .A2(n1683), .A3(
        write_data[23]), .A4(n3056), .Y(\words[25]/data_i[23] ) );
  AO22X1_RVT U4573 ( .A1(\read_value_mux[25][24] ), .A2(n1683), .A3(
        write_data[24]), .A4(n3056), .Y(\words[25]/data_i[24] ) );
  AO22X1_RVT U4574 ( .A1(\read_value_mux[25][25] ), .A2(n1683), .A3(
        write_data[25]), .A4(n3056), .Y(\words[25]/data_i[25] ) );
  AO22X1_RVT U4575 ( .A1(\read_value_mux[25][26] ), .A2(n1683), .A3(
        write_data[26]), .A4(n3056), .Y(\words[25]/data_i[26] ) );
  AO22X1_RVT U4576 ( .A1(\read_value_mux[25][27] ), .A2(n1683), .A3(
        write_data[27]), .A4(n3056), .Y(\words[25]/data_i[27] ) );
  AO22X1_RVT U4577 ( .A1(\read_value_mux[25][28] ), .A2(n1683), .A3(
        write_data[28]), .A4(n3056), .Y(\words[25]/data_i[28] ) );
  AO22X1_RVT U4578 ( .A1(\read_value_mux[25][29] ), .A2(n1683), .A3(
        write_data[29]), .A4(n3056), .Y(\words[25]/data_i[29] ) );
  AO22X1_RVT U4579 ( .A1(\read_value_mux[25][2] ), .A2(n1683), .A3(
        write_data[2]), .A4(n3056), .Y(\words[25]/data_i[2] ) );
  AO22X1_RVT U4580 ( .A1(n3056), .A2(write_data[30]), .A3(
        \read_value_mux[25][30] ), .A4(n1683), .Y(\words[25]/data_i[30] ) );
  AO22X1_RVT U4581 ( .A1(\read_value_mux[25][31] ), .A2(n1683), .A3(
        write_data[31]), .A4(n3056), .Y(\words[25]/data_i[31] ) );
  AO22X1_RVT U4582 ( .A1(\read_value_mux[25][3] ), .A2(n1683), .A3(
        write_data[3]), .A4(n3056), .Y(\words[25]/data_i[3] ) );
  AO22X1_RVT U4583 ( .A1(\read_value_mux[25][4] ), .A2(n1683), .A3(
        write_data[4]), .A4(n3056), .Y(\words[25]/data_i[4] ) );
  AO22X1_RVT U4584 ( .A1(\read_value_mux[25][5] ), .A2(n1683), .A3(
        write_data[5]), .A4(n3056), .Y(\words[25]/data_i[5] ) );
  AO22X1_RVT U4585 ( .A1(\read_value_mux[25][6] ), .A2(n1683), .A3(
        write_data[6]), .A4(n3056), .Y(\words[25]/data_i[6] ) );
  AO22X1_RVT U4586 ( .A1(\read_value_mux[25][7] ), .A2(n1683), .A3(
        write_data[7]), .A4(n3056), .Y(\words[25]/data_i[7] ) );
  AO22X1_RVT U4587 ( .A1(\read_value_mux[25][8] ), .A2(n1683), .A3(
        write_data[8]), .A4(n3056), .Y(\words[25]/data_i[8] ) );
  AO22X1_RVT U4588 ( .A1(\read_value_mux[25][9] ), .A2(n1683), .A3(
        write_data[9]), .A4(n3056), .Y(\words[25]/data_i[9] ) );
  AO21X1_RVT U4589 ( .A1(\words[25]/valid_o ), .A2(n1683), .A3(n3056), .Y(
        \words[25]/valid_i ) );
  AO22X1_RVT U4590 ( .A1(\read_value_mux[26][0] ), .A2(n3058), .A3(
        write_data[0]), .A4(n3057), .Y(\words[26]/data_i[0] ) );
  AO22X1_RVT U4591 ( .A1(\read_value_mux[26][10] ), .A2(n3058), .A3(
        write_data[10]), .A4(n3057), .Y(\words[26]/data_i[10] ) );
  AO22X1_RVT U4592 ( .A1(\read_value_mux[26][11] ), .A2(n3058), .A3(
        write_data[11]), .A4(n3057), .Y(\words[26]/data_i[11] ) );
  AO22X1_RVT U4593 ( .A1(\read_value_mux[26][12] ), .A2(n3058), .A3(
        write_data[12]), .A4(n3057), .Y(\words[26]/data_i[12] ) );
  AO22X1_RVT U4594 ( .A1(\read_value_mux[26][13] ), .A2(n3058), .A3(
        write_data[13]), .A4(n3057), .Y(\words[26]/data_i[13] ) );
  AO22X1_RVT U4595 ( .A1(\read_value_mux[26][14] ), .A2(n3058), .A3(
        write_data[14]), .A4(n3057), .Y(\words[26]/data_i[14] ) );
  AO22X1_RVT U4596 ( .A1(\read_value_mux[26][15] ), .A2(n3058), .A3(
        write_data[15]), .A4(n3057), .Y(\words[26]/data_i[15] ) );
  AO22X1_RVT U4597 ( .A1(\read_value_mux[26][16] ), .A2(n3058), .A3(
        write_data[16]), .A4(n3057), .Y(\words[26]/data_i[16] ) );
  AO22X1_RVT U4598 ( .A1(\read_value_mux[26][17] ), .A2(n3058), .A3(
        write_data[17]), .A4(n3057), .Y(\words[26]/data_i[17] ) );
  AO22X1_RVT U4599 ( .A1(\read_value_mux[26][18] ), .A2(n3058), .A3(
        write_data[18]), .A4(n3057), .Y(\words[26]/data_i[18] ) );
  AO22X1_RVT U4600 ( .A1(\read_value_mux[26][19] ), .A2(n3058), .A3(
        write_data[19]), .A4(n3057), .Y(\words[26]/data_i[19] ) );
  AO22X1_RVT U4601 ( .A1(n3057), .A2(write_data[1]), .A3(
        \read_value_mux[26][1] ), .A4(n3058), .Y(\words[26]/data_i[1] ) );
  AO22X1_RVT U4602 ( .A1(\read_value_mux[26][20] ), .A2(n3058), .A3(
        write_data[20]), .A4(n3057), .Y(\words[26]/data_i[20] ) );
  AO22X1_RVT U4603 ( .A1(\read_value_mux[26][21] ), .A2(n3058), .A3(
        write_data[21]), .A4(n3057), .Y(\words[26]/data_i[21] ) );
  AO22X1_RVT U4604 ( .A1(\read_value_mux[26][22] ), .A2(n3058), .A3(
        write_data[22]), .A4(n3057), .Y(\words[26]/data_i[22] ) );
  AO22X1_RVT U4605 ( .A1(\read_value_mux[26][23] ), .A2(n3058), .A3(
        write_data[23]), .A4(n3057), .Y(\words[26]/data_i[23] ) );
  AO22X1_RVT U4606 ( .A1(\read_value_mux[26][24] ), .A2(n3058), .A3(
        write_data[24]), .A4(n3057), .Y(\words[26]/data_i[24] ) );
  AO22X1_RVT U4607 ( .A1(\read_value_mux[26][25] ), .A2(n3058), .A3(
        write_data[25]), .A4(n3057), .Y(\words[26]/data_i[25] ) );
  AO22X1_RVT U4608 ( .A1(\read_value_mux[26][26] ), .A2(n3058), .A3(
        write_data[26]), .A4(n3057), .Y(\words[26]/data_i[26] ) );
  AO22X1_RVT U4609 ( .A1(\read_value_mux[26][27] ), .A2(n3058), .A3(
        write_data[27]), .A4(n3057), .Y(\words[26]/data_i[27] ) );
  AO22X1_RVT U4610 ( .A1(\read_value_mux[26][28] ), .A2(n3058), .A3(
        write_data[28]), .A4(n3057), .Y(\words[26]/data_i[28] ) );
  AO22X1_RVT U4611 ( .A1(\read_value_mux[26][29] ), .A2(n3058), .A3(
        write_data[29]), .A4(n3057), .Y(\words[26]/data_i[29] ) );
  AO22X1_RVT U4612 ( .A1(\read_value_mux[26][2] ), .A2(n3058), .A3(
        write_data[2]), .A4(n3057), .Y(\words[26]/data_i[2] ) );
  AO22X1_RVT U4613 ( .A1(n3057), .A2(write_data[30]), .A3(
        \read_value_mux[26][30] ), .A4(n3058), .Y(\words[26]/data_i[30] ) );
  AO22X1_RVT U4614 ( .A1(\read_value_mux[26][31] ), .A2(n3058), .A3(
        write_data[31]), .A4(n3057), .Y(\words[26]/data_i[31] ) );
  AO22X1_RVT U4615 ( .A1(\read_value_mux[26][3] ), .A2(n3058), .A3(
        write_data[3]), .A4(n3057), .Y(\words[26]/data_i[3] ) );
  AO22X1_RVT U4616 ( .A1(\read_value_mux[26][4] ), .A2(n3058), .A3(
        write_data[4]), .A4(n3057), .Y(\words[26]/data_i[4] ) );
  AO22X1_RVT U4617 ( .A1(\read_value_mux[26][5] ), .A2(n3058), .A3(
        write_data[5]), .A4(n3057), .Y(\words[26]/data_i[5] ) );
  AO22X1_RVT U4618 ( .A1(\read_value_mux[26][6] ), .A2(n3058), .A3(
        write_data[6]), .A4(n3057), .Y(\words[26]/data_i[6] ) );
  AO22X1_RVT U4619 ( .A1(\read_value_mux[26][7] ), .A2(n3058), .A3(
        write_data[7]), .A4(n3057), .Y(\words[26]/data_i[7] ) );
  AO22X1_RVT U4620 ( .A1(\read_value_mux[26][8] ), .A2(n3058), .A3(
        write_data[8]), .A4(n3057), .Y(\words[26]/data_i[8] ) );
  AO22X1_RVT U4621 ( .A1(\read_value_mux[26][9] ), .A2(n3058), .A3(
        write_data[9]), .A4(n3057), .Y(\words[26]/data_i[9] ) );
  AO21X1_RVT U4622 ( .A1(\words[26]/valid_o ), .A2(n3058), .A3(n3057), .Y(
        \words[26]/valid_i ) );
  AO22X1_RVT U4623 ( .A1(\read_value_mux[27][0] ), .A2(n1633), .A3(
        write_data[0]), .A4(n3061), .Y(\words[27]/data_i[0] ) );
  AO22X1_RVT U4624 ( .A1(\read_value_mux[27][10] ), .A2(n1633), .A3(
        write_data[10]), .A4(n3061), .Y(\words[27]/data_i[10] ) );
  AO22X1_RVT U4625 ( .A1(\read_value_mux[27][11] ), .A2(n1633), .A3(
        write_data[11]), .A4(n3061), .Y(\words[27]/data_i[11] ) );
  AO22X1_RVT U4626 ( .A1(\read_value_mux[27][12] ), .A2(n1633), .A3(
        write_data[12]), .A4(n3061), .Y(\words[27]/data_i[12] ) );
  AO22X1_RVT U4627 ( .A1(\read_value_mux[27][13] ), .A2(n1633), .A3(
        write_data[13]), .A4(n3061), .Y(\words[27]/data_i[13] ) );
  AO22X1_RVT U4628 ( .A1(\read_value_mux[27][14] ), .A2(n1633), .A3(
        write_data[14]), .A4(n3061), .Y(\words[27]/data_i[14] ) );
  AO22X1_RVT U4629 ( .A1(\read_value_mux[27][15] ), .A2(n1633), .A3(
        write_data[15]), .A4(n3061), .Y(\words[27]/data_i[15] ) );
  AO22X1_RVT U4630 ( .A1(\read_value_mux[27][16] ), .A2(n1633), .A3(
        write_data[16]), .A4(n3061), .Y(\words[27]/data_i[16] ) );
  AO22X1_RVT U4631 ( .A1(\read_value_mux[27][17] ), .A2(n1633), .A3(
        write_data[17]), .A4(n3061), .Y(\words[27]/data_i[17] ) );
  AO22X1_RVT U4632 ( .A1(\read_value_mux[27][18] ), .A2(n1633), .A3(
        write_data[18]), .A4(n3061), .Y(\words[27]/data_i[18] ) );
  AO22X1_RVT U4633 ( .A1(\read_value_mux[27][19] ), .A2(n1633), .A3(
        write_data[19]), .A4(n3061), .Y(\words[27]/data_i[19] ) );
  AO22X1_RVT U4634 ( .A1(n3061), .A2(write_data[1]), .A3(
        \read_value_mux[27][1] ), .A4(n1633), .Y(\words[27]/data_i[1] ) );
  AO22X1_RVT U4635 ( .A1(\read_value_mux[27][20] ), .A2(n1633), .A3(
        write_data[20]), .A4(n3061), .Y(\words[27]/data_i[20] ) );
  AO22X1_RVT U4636 ( .A1(\read_value_mux[27][21] ), .A2(n1633), .A3(
        write_data[21]), .A4(n3061), .Y(\words[27]/data_i[21] ) );
  AO22X1_RVT U4637 ( .A1(\read_value_mux[27][22] ), .A2(n1633), .A3(
        write_data[22]), .A4(n3061), .Y(\words[27]/data_i[22] ) );
  AO22X1_RVT U4638 ( .A1(\read_value_mux[27][23] ), .A2(n1633), .A3(
        write_data[23]), .A4(n3061), .Y(\words[27]/data_i[23] ) );
  AO22X1_RVT U4639 ( .A1(\read_value_mux[27][24] ), .A2(n1633), .A3(
        write_data[24]), .A4(n3061), .Y(\words[27]/data_i[24] ) );
  AO22X1_RVT U4640 ( .A1(\read_value_mux[27][25] ), .A2(n1633), .A3(
        write_data[25]), .A4(n3061), .Y(\words[27]/data_i[25] ) );
  AO22X1_RVT U4641 ( .A1(\read_value_mux[27][26] ), .A2(n1633), .A3(
        write_data[26]), .A4(n3061), .Y(\words[27]/data_i[26] ) );
  AO22X1_RVT U4642 ( .A1(\read_value_mux[27][27] ), .A2(n1633), .A3(
        write_data[27]), .A4(n3061), .Y(\words[27]/data_i[27] ) );
  AO22X1_RVT U4643 ( .A1(\read_value_mux[27][28] ), .A2(n1633), .A3(
        write_data[28]), .A4(n3061), .Y(\words[27]/data_i[28] ) );
  AO22X1_RVT U4644 ( .A1(\read_value_mux[27][29] ), .A2(n1633), .A3(
        write_data[29]), .A4(n3061), .Y(\words[27]/data_i[29] ) );
  AO22X1_RVT U4645 ( .A1(\read_value_mux[27][2] ), .A2(n1633), .A3(
        write_data[2]), .A4(n3061), .Y(\words[27]/data_i[2] ) );
  AO22X1_RVT U4646 ( .A1(n3061), .A2(write_data[30]), .A3(
        \read_value_mux[27][30] ), .A4(n1633), .Y(\words[27]/data_i[30] ) );
  AO22X1_RVT U4647 ( .A1(\read_value_mux[27][31] ), .A2(n1633), .A3(
        write_data[31]), .A4(n3061), .Y(\words[27]/data_i[31] ) );
  AO22X1_RVT U4648 ( .A1(\read_value_mux[27][3] ), .A2(n1633), .A3(
        write_data[3]), .A4(n3061), .Y(\words[27]/data_i[3] ) );
  AO22X1_RVT U4649 ( .A1(\read_value_mux[27][4] ), .A2(n1633), .A3(
        write_data[4]), .A4(n3061), .Y(\words[27]/data_i[4] ) );
  AO22X1_RVT U4650 ( .A1(\read_value_mux[27][5] ), .A2(n1633), .A3(
        write_data[5]), .A4(n3061), .Y(\words[27]/data_i[5] ) );
  AO22X1_RVT U4651 ( .A1(\read_value_mux[27][6] ), .A2(n1633), .A3(
        write_data[6]), .A4(n3061), .Y(\words[27]/data_i[6] ) );
  AO22X1_RVT U4652 ( .A1(\read_value_mux[27][7] ), .A2(n1633), .A3(
        write_data[7]), .A4(n3061), .Y(\words[27]/data_i[7] ) );
  AO22X1_RVT U4653 ( .A1(\read_value_mux[27][8] ), .A2(n1633), .A3(
        write_data[8]), .A4(n3061), .Y(\words[27]/data_i[8] ) );
  AO22X1_RVT U4654 ( .A1(\read_value_mux[27][9] ), .A2(n1633), .A3(
        write_data[9]), .A4(n3061), .Y(\words[27]/data_i[9] ) );
  AO21X1_RVT U4655 ( .A1(\words[27]/valid_o ), .A2(n1633), .A3(n3061), .Y(
        \words[27]/valid_i ) );
  AO22X1_RVT U4656 ( .A1(\read_value_mux[28][0] ), .A2(n1678), .A3(
        write_data[0]), .A4(n3062), .Y(\words[28]/data_i[0] ) );
  AO22X1_RVT U4657 ( .A1(\read_value_mux[28][10] ), .A2(n1678), .A3(
        write_data[10]), .A4(n3062), .Y(\words[28]/data_i[10] ) );
  AO22X1_RVT U4658 ( .A1(\read_value_mux[28][11] ), .A2(n1678), .A3(
        write_data[11]), .A4(n3062), .Y(\words[28]/data_i[11] ) );
  AO22X1_RVT U4659 ( .A1(\read_value_mux[28][12] ), .A2(n1678), .A3(
        write_data[12]), .A4(n3062), .Y(\words[28]/data_i[12] ) );
  AO22X1_RVT U4660 ( .A1(\read_value_mux[28][13] ), .A2(n1678), .A3(
        write_data[13]), .A4(n3062), .Y(\words[28]/data_i[13] ) );
  AO22X1_RVT U4661 ( .A1(\read_value_mux[28][14] ), .A2(n1678), .A3(
        write_data[14]), .A4(n3062), .Y(\words[28]/data_i[14] ) );
  AO22X1_RVT U4662 ( .A1(\read_value_mux[28][15] ), .A2(n1678), .A3(
        write_data[15]), .A4(n3062), .Y(\words[28]/data_i[15] ) );
  AO22X1_RVT U4663 ( .A1(\read_value_mux[28][16] ), .A2(n1678), .A3(
        write_data[16]), .A4(n3062), .Y(\words[28]/data_i[16] ) );
  AO22X1_RVT U4664 ( .A1(\read_value_mux[28][17] ), .A2(n1678), .A3(
        write_data[17]), .A4(n3062), .Y(\words[28]/data_i[17] ) );
  AO22X1_RVT U4665 ( .A1(\read_value_mux[28][18] ), .A2(n1678), .A3(
        write_data[18]), .A4(n3062), .Y(\words[28]/data_i[18] ) );
  AO22X1_RVT U4666 ( .A1(\read_value_mux[28][19] ), .A2(n1678), .A3(
        write_data[19]), .A4(n3062), .Y(\words[28]/data_i[19] ) );
  AO22X1_RVT U4667 ( .A1(n3062), .A2(write_data[1]), .A3(
        \read_value_mux[28][1] ), .A4(n1678), .Y(\words[28]/data_i[1] ) );
  AO22X1_RVT U4668 ( .A1(\read_value_mux[28][20] ), .A2(n1678), .A3(
        write_data[20]), .A4(n3062), .Y(\words[28]/data_i[20] ) );
  AO22X1_RVT U4669 ( .A1(\read_value_mux[28][21] ), .A2(n1678), .A3(
        write_data[21]), .A4(n3062), .Y(\words[28]/data_i[21] ) );
  AO22X1_RVT U4670 ( .A1(\read_value_mux[28][22] ), .A2(n1678), .A3(
        write_data[22]), .A4(n3062), .Y(\words[28]/data_i[22] ) );
  AO22X1_RVT U4671 ( .A1(\read_value_mux[28][23] ), .A2(n1678), .A3(
        write_data[23]), .A4(n3062), .Y(\words[28]/data_i[23] ) );
  AO22X1_RVT U4672 ( .A1(\read_value_mux[28][24] ), .A2(n1678), .A3(
        write_data[24]), .A4(n3062), .Y(\words[28]/data_i[24] ) );
  AO22X1_RVT U4673 ( .A1(\read_value_mux[28][25] ), .A2(n1678), .A3(
        write_data[25]), .A4(n3062), .Y(\words[28]/data_i[25] ) );
  AO22X1_RVT U4674 ( .A1(\read_value_mux[28][26] ), .A2(n1678), .A3(
        write_data[26]), .A4(n3062), .Y(\words[28]/data_i[26] ) );
  AO22X1_RVT U4675 ( .A1(\read_value_mux[28][27] ), .A2(n1678), .A3(
        write_data[27]), .A4(n3062), .Y(\words[28]/data_i[27] ) );
  AO22X1_RVT U4676 ( .A1(\read_value_mux[28][28] ), .A2(n1678), .A3(
        write_data[28]), .A4(n3062), .Y(\words[28]/data_i[28] ) );
  AO22X1_RVT U4677 ( .A1(\read_value_mux[28][29] ), .A2(n1678), .A3(
        write_data[29]), .A4(n3062), .Y(\words[28]/data_i[29] ) );
  AO22X1_RVT U4678 ( .A1(\read_value_mux[28][2] ), .A2(n1678), .A3(
        write_data[2]), .A4(n3062), .Y(\words[28]/data_i[2] ) );
  AO22X1_RVT U4679 ( .A1(n3062), .A2(write_data[30]), .A3(
        \read_value_mux[28][30] ), .A4(n1678), .Y(\words[28]/data_i[30] ) );
  AO22X1_RVT U4680 ( .A1(\read_value_mux[28][31] ), .A2(n1678), .A3(
        write_data[31]), .A4(n3062), .Y(\words[28]/data_i[31] ) );
  AO22X1_RVT U4681 ( .A1(\read_value_mux[28][3] ), .A2(n1678), .A3(
        write_data[3]), .A4(n3062), .Y(\words[28]/data_i[3] ) );
  AO22X1_RVT U4682 ( .A1(\read_value_mux[28][4] ), .A2(n1678), .A3(
        write_data[4]), .A4(n3062), .Y(\words[28]/data_i[4] ) );
  AO22X1_RVT U4683 ( .A1(\read_value_mux[28][5] ), .A2(n1678), .A3(
        write_data[5]), .A4(n3062), .Y(\words[28]/data_i[5] ) );
  AO22X1_RVT U4684 ( .A1(\read_value_mux[28][6] ), .A2(n1678), .A3(
        write_data[6]), .A4(n3062), .Y(\words[28]/data_i[6] ) );
  AO22X1_RVT U4685 ( .A1(\read_value_mux[28][7] ), .A2(n1678), .A3(
        write_data[7]), .A4(n3062), .Y(\words[28]/data_i[7] ) );
  AO22X1_RVT U4686 ( .A1(\read_value_mux[28][8] ), .A2(n1678), .A3(
        write_data[8]), .A4(n3062), .Y(\words[28]/data_i[8] ) );
  AO22X1_RVT U4687 ( .A1(\read_value_mux[28][9] ), .A2(n1678), .A3(
        write_data[9]), .A4(n3062), .Y(\words[28]/data_i[9] ) );
  AO21X1_RVT U4688 ( .A1(\words[28]/valid_o ), .A2(n1678), .A3(n3062), .Y(
        \words[28]/valid_i ) );
  AO22X1_RVT U4689 ( .A1(\read_value_mux[29][0] ), .A2(n3064), .A3(
        write_data[0]), .A4(n3063), .Y(\words[29]/data_i[0] ) );
  AO22X1_RVT U4690 ( .A1(\read_value_mux[29][10] ), .A2(n3064), .A3(
        write_data[10]), .A4(n3063), .Y(\words[29]/data_i[10] ) );
  AO22X1_RVT U4691 ( .A1(\read_value_mux[29][11] ), .A2(n3064), .A3(
        write_data[11]), .A4(n3063), .Y(\words[29]/data_i[11] ) );
  AO22X1_RVT U4692 ( .A1(\read_value_mux[29][12] ), .A2(n3064), .A3(
        write_data[12]), .A4(n3063), .Y(\words[29]/data_i[12] ) );
  AO22X1_RVT U4693 ( .A1(\read_value_mux[29][13] ), .A2(n3064), .A3(
        write_data[13]), .A4(n3063), .Y(\words[29]/data_i[13] ) );
  AO22X1_RVT U4694 ( .A1(\read_value_mux[29][14] ), .A2(n3064), .A3(
        write_data[14]), .A4(n3063), .Y(\words[29]/data_i[14] ) );
  AO22X1_RVT U4695 ( .A1(\read_value_mux[29][15] ), .A2(n3064), .A3(
        write_data[15]), .A4(n3063), .Y(\words[29]/data_i[15] ) );
  AO22X1_RVT U4696 ( .A1(\read_value_mux[29][16] ), .A2(n3064), .A3(
        write_data[16]), .A4(n3063), .Y(\words[29]/data_i[16] ) );
  AO22X1_RVT U4697 ( .A1(\read_value_mux[29][17] ), .A2(n3064), .A3(
        write_data[17]), .A4(n3063), .Y(\words[29]/data_i[17] ) );
  AO22X1_RVT U4698 ( .A1(\read_value_mux[29][18] ), .A2(n3064), .A3(
        write_data[18]), .A4(n3063), .Y(\words[29]/data_i[18] ) );
  AO22X1_RVT U4699 ( .A1(\read_value_mux[29][19] ), .A2(n3064), .A3(
        write_data[19]), .A4(n3063), .Y(\words[29]/data_i[19] ) );
  AO22X1_RVT U4700 ( .A1(n3063), .A2(write_data[1]), .A3(
        \read_value_mux[29][1] ), .A4(n3064), .Y(\words[29]/data_i[1] ) );
  AO22X1_RVT U4701 ( .A1(\read_value_mux[29][20] ), .A2(n3064), .A3(
        write_data[20]), .A4(n3063), .Y(\words[29]/data_i[20] ) );
  AO22X1_RVT U4702 ( .A1(\read_value_mux[29][21] ), .A2(n3064), .A3(
        write_data[21]), .A4(n3063), .Y(\words[29]/data_i[21] ) );
  AO22X1_RVT U4703 ( .A1(\read_value_mux[29][22] ), .A2(n3064), .A3(
        write_data[22]), .A4(n3063), .Y(\words[29]/data_i[22] ) );
  AO22X1_RVT U4704 ( .A1(\read_value_mux[29][23] ), .A2(n3064), .A3(
        write_data[23]), .A4(n3063), .Y(\words[29]/data_i[23] ) );
  AO22X1_RVT U4705 ( .A1(\read_value_mux[29][24] ), .A2(n3064), .A3(
        write_data[24]), .A4(n3063), .Y(\words[29]/data_i[24] ) );
  AO22X1_RVT U4706 ( .A1(\read_value_mux[29][25] ), .A2(n3064), .A3(
        write_data[25]), .A4(n3063), .Y(\words[29]/data_i[25] ) );
  AO22X1_RVT U4707 ( .A1(\read_value_mux[29][26] ), .A2(n3064), .A3(
        write_data[26]), .A4(n3063), .Y(\words[29]/data_i[26] ) );
  AO22X1_RVT U4708 ( .A1(\read_value_mux[29][27] ), .A2(n3064), .A3(
        write_data[27]), .A4(n3063), .Y(\words[29]/data_i[27] ) );
  AO22X1_RVT U4709 ( .A1(\read_value_mux[29][28] ), .A2(n3064), .A3(
        write_data[28]), .A4(n3063), .Y(\words[29]/data_i[28] ) );
  AO22X1_RVT U4710 ( .A1(\read_value_mux[29][29] ), .A2(n3064), .A3(
        write_data[29]), .A4(n3063), .Y(\words[29]/data_i[29] ) );
  AO22X1_RVT U4711 ( .A1(\read_value_mux[29][2] ), .A2(n3064), .A3(
        write_data[2]), .A4(n3063), .Y(\words[29]/data_i[2] ) );
  AO22X1_RVT U4712 ( .A1(n3063), .A2(write_data[30]), .A3(
        \read_value_mux[29][30] ), .A4(n3064), .Y(\words[29]/data_i[30] ) );
  AO22X1_RVT U4713 ( .A1(\read_value_mux[29][31] ), .A2(n3064), .A3(
        write_data[31]), .A4(n3063), .Y(\words[29]/data_i[31] ) );
  AO22X1_RVT U4714 ( .A1(\read_value_mux[29][3] ), .A2(n3064), .A3(
        write_data[3]), .A4(n3063), .Y(\words[29]/data_i[3] ) );
  AO22X1_RVT U4715 ( .A1(\read_value_mux[29][4] ), .A2(n3064), .A3(
        write_data[4]), .A4(n3063), .Y(\words[29]/data_i[4] ) );
  AO22X1_RVT U4716 ( .A1(\read_value_mux[29][5] ), .A2(n3064), .A3(
        write_data[5]), .A4(n3063), .Y(\words[29]/data_i[5] ) );
  AO22X1_RVT U4717 ( .A1(\read_value_mux[29][6] ), .A2(n3064), .A3(
        write_data[6]), .A4(n3063), .Y(\words[29]/data_i[6] ) );
  AO22X1_RVT U4718 ( .A1(\read_value_mux[29][7] ), .A2(n3064), .A3(
        write_data[7]), .A4(n3063), .Y(\words[29]/data_i[7] ) );
  AO22X1_RVT U4719 ( .A1(\read_value_mux[29][8] ), .A2(n3064), .A3(
        write_data[8]), .A4(n3063), .Y(\words[29]/data_i[8] ) );
  AO22X1_RVT U4720 ( .A1(\read_value_mux[29][9] ), .A2(n3064), .A3(
        write_data[9]), .A4(n3063), .Y(\words[29]/data_i[9] ) );
  AO21X1_RVT U4721 ( .A1(\words[29]/valid_o ), .A2(n3064), .A3(n3063), .Y(
        \words[29]/valid_i ) );
  AO22X1_RVT U4722 ( .A1(\read_value_mux[2][0] ), .A2(n1687), .A3(
        write_data[0]), .A4(n3065), .Y(\words[2]/data_i[0] ) );
  AO22X1_RVT U4723 ( .A1(\read_value_mux[2][10] ), .A2(n1687), .A3(
        write_data[10]), .A4(n3065), .Y(\words[2]/data_i[10] ) );
  AO22X1_RVT U4724 ( .A1(\read_value_mux[2][11] ), .A2(n1687), .A3(
        write_data[11]), .A4(n3065), .Y(\words[2]/data_i[11] ) );
  AO22X1_RVT U4725 ( .A1(\read_value_mux[2][12] ), .A2(n1687), .A3(
        write_data[12]), .A4(n3065), .Y(\words[2]/data_i[12] ) );
  AO22X1_RVT U4726 ( .A1(\read_value_mux[2][13] ), .A2(n1687), .A3(
        write_data[13]), .A4(n3065), .Y(\words[2]/data_i[13] ) );
  AO22X1_RVT U4727 ( .A1(\read_value_mux[2][14] ), .A2(n1687), .A3(
        write_data[14]), .A4(n3065), .Y(\words[2]/data_i[14] ) );
  AO22X1_RVT U4728 ( .A1(\read_value_mux[2][15] ), .A2(n1687), .A3(
        write_data[15]), .A4(n3065), .Y(\words[2]/data_i[15] ) );
  AO22X1_RVT U4729 ( .A1(\read_value_mux[2][16] ), .A2(n1687), .A3(
        write_data[16]), .A4(n3065), .Y(\words[2]/data_i[16] ) );
  AO22X1_RVT U4730 ( .A1(\read_value_mux[2][17] ), .A2(n1687), .A3(
        write_data[17]), .A4(n3065), .Y(\words[2]/data_i[17] ) );
  AO22X1_RVT U4731 ( .A1(\read_value_mux[2][18] ), .A2(n1687), .A3(
        write_data[18]), .A4(n3065), .Y(\words[2]/data_i[18] ) );
  AO22X1_RVT U4732 ( .A1(\read_value_mux[2][19] ), .A2(n1687), .A3(
        write_data[19]), .A4(n3065), .Y(\words[2]/data_i[19] ) );
  AO22X1_RVT U4733 ( .A1(n3065), .A2(write_data[1]), .A3(
        \read_value_mux[2][1] ), .A4(n1687), .Y(\words[2]/data_i[1] ) );
  AO22X1_RVT U4734 ( .A1(\read_value_mux[2][20] ), .A2(n1687), .A3(
        write_data[20]), .A4(n3065), .Y(\words[2]/data_i[20] ) );
  AO22X1_RVT U4735 ( .A1(\read_value_mux[2][21] ), .A2(n1687), .A3(
        write_data[21]), .A4(n3065), .Y(\words[2]/data_i[21] ) );
  AO22X1_RVT U4736 ( .A1(\read_value_mux[2][22] ), .A2(n1687), .A3(
        write_data[22]), .A4(n3065), .Y(\words[2]/data_i[22] ) );
  AO22X1_RVT U4737 ( .A1(\read_value_mux[2][23] ), .A2(n1687), .A3(
        write_data[23]), .A4(n3065), .Y(\words[2]/data_i[23] ) );
  AO22X1_RVT U4738 ( .A1(\read_value_mux[2][24] ), .A2(n1687), .A3(
        write_data[24]), .A4(n3065), .Y(\words[2]/data_i[24] ) );
  AO22X1_RVT U4739 ( .A1(\read_value_mux[2][25] ), .A2(n1687), .A3(
        write_data[25]), .A4(n3065), .Y(\words[2]/data_i[25] ) );
  AO22X1_RVT U4740 ( .A1(\read_value_mux[2][26] ), .A2(n1687), .A3(
        write_data[26]), .A4(n3065), .Y(\words[2]/data_i[26] ) );
  AO22X1_RVT U4741 ( .A1(\read_value_mux[2][27] ), .A2(n1687), .A3(
        write_data[27]), .A4(n3065), .Y(\words[2]/data_i[27] ) );
  AO22X1_RVT U4742 ( .A1(\read_value_mux[2][28] ), .A2(n1687), .A3(
        write_data[28]), .A4(n3065), .Y(\words[2]/data_i[28] ) );
  AO22X1_RVT U4743 ( .A1(\read_value_mux[2][29] ), .A2(n1687), .A3(
        write_data[29]), .A4(n3065), .Y(\words[2]/data_i[29] ) );
  AO22X1_RVT U4744 ( .A1(\read_value_mux[2][2] ), .A2(n1687), .A3(
        write_data[2]), .A4(n3065), .Y(\words[2]/data_i[2] ) );
  AO22X1_RVT U4745 ( .A1(n3065), .A2(write_data[30]), .A3(
        \read_value_mux[2][30] ), .A4(n1687), .Y(\words[2]/data_i[30] ) );
  AO22X1_RVT U4746 ( .A1(\read_value_mux[2][31] ), .A2(n1687), .A3(
        write_data[31]), .A4(n3065), .Y(\words[2]/data_i[31] ) );
  AO22X1_RVT U4747 ( .A1(\read_value_mux[2][3] ), .A2(n1687), .A3(
        write_data[3]), .A4(n3065), .Y(\words[2]/data_i[3] ) );
  AO22X1_RVT U4748 ( .A1(\read_value_mux[2][4] ), .A2(n1687), .A3(
        write_data[4]), .A4(n3065), .Y(\words[2]/data_i[4] ) );
  AO22X1_RVT U4749 ( .A1(\read_value_mux[2][5] ), .A2(n1687), .A3(
        write_data[5]), .A4(n3065), .Y(\words[2]/data_i[5] ) );
  AO22X1_RVT U4750 ( .A1(\read_value_mux[2][6] ), .A2(n1687), .A3(
        write_data[6]), .A4(n3065), .Y(\words[2]/data_i[6] ) );
  AO22X1_RVT U4751 ( .A1(\read_value_mux[2][7] ), .A2(n1687), .A3(
        write_data[7]), .A4(n3065), .Y(\words[2]/data_i[7] ) );
  AO22X1_RVT U4752 ( .A1(\read_value_mux[2][8] ), .A2(n1687), .A3(
        write_data[8]), .A4(n3065), .Y(\words[2]/data_i[8] ) );
  AO22X1_RVT U4753 ( .A1(\read_value_mux[2][9] ), .A2(n1687), .A3(
        write_data[9]), .A4(n3065), .Y(\words[2]/data_i[9] ) );
  AO21X1_RVT U4754 ( .A1(\words[2]/valid_o ), .A2(n1687), .A3(n3065), .Y(
        \words[2]/valid_i ) );
  AO22X1_RVT U4755 ( .A1(\read_value_mux[30][0] ), .A2(n3067), .A3(
        write_data[0]), .A4(n3066), .Y(\words[30]/data_i[0] ) );
  AO22X1_RVT U4756 ( .A1(\read_value_mux[30][10] ), .A2(n3067), .A3(
        write_data[10]), .A4(n3066), .Y(\words[30]/data_i[10] ) );
  AO22X1_RVT U4757 ( .A1(\read_value_mux[30][11] ), .A2(n3067), .A3(
        write_data[11]), .A4(n3066), .Y(\words[30]/data_i[11] ) );
  AO22X1_RVT U4758 ( .A1(\read_value_mux[30][12] ), .A2(n3067), .A3(
        write_data[12]), .A4(n3066), .Y(\words[30]/data_i[12] ) );
  AO22X1_RVT U4759 ( .A1(\read_value_mux[30][13] ), .A2(n3067), .A3(
        write_data[13]), .A4(n3066), .Y(\words[30]/data_i[13] ) );
  AO22X1_RVT U4760 ( .A1(\read_value_mux[30][14] ), .A2(n3067), .A3(
        write_data[14]), .A4(n3066), .Y(\words[30]/data_i[14] ) );
  AO22X1_RVT U4761 ( .A1(\read_value_mux[30][15] ), .A2(n3067), .A3(
        write_data[15]), .A4(n3066), .Y(\words[30]/data_i[15] ) );
  AO22X1_RVT U4762 ( .A1(\read_value_mux[30][16] ), .A2(n3067), .A3(
        write_data[16]), .A4(n3066), .Y(\words[30]/data_i[16] ) );
  AO22X1_RVT U4763 ( .A1(\read_value_mux[30][17] ), .A2(n3067), .A3(
        write_data[17]), .A4(n3066), .Y(\words[30]/data_i[17] ) );
  AO22X1_RVT U4764 ( .A1(\read_value_mux[30][18] ), .A2(n3067), .A3(
        write_data[18]), .A4(n3066), .Y(\words[30]/data_i[18] ) );
  AO22X1_RVT U4765 ( .A1(\read_value_mux[30][19] ), .A2(n3067), .A3(
        write_data[19]), .A4(n3066), .Y(\words[30]/data_i[19] ) );
  AO22X1_RVT U4766 ( .A1(n3066), .A2(write_data[1]), .A3(
        \read_value_mux[30][1] ), .A4(n3067), .Y(\words[30]/data_i[1] ) );
  AO22X1_RVT U4767 ( .A1(\read_value_mux[30][20] ), .A2(n3067), .A3(
        write_data[20]), .A4(n3066), .Y(\words[30]/data_i[20] ) );
  AO22X1_RVT U4768 ( .A1(\read_value_mux[30][21] ), .A2(n3067), .A3(
        write_data[21]), .A4(n3066), .Y(\words[30]/data_i[21] ) );
  AO22X1_RVT U4769 ( .A1(\read_value_mux[30][22] ), .A2(n3067), .A3(
        write_data[22]), .A4(n3066), .Y(\words[30]/data_i[22] ) );
  AO22X1_RVT U4770 ( .A1(\read_value_mux[30][23] ), .A2(n3067), .A3(
        write_data[23]), .A4(n3066), .Y(\words[30]/data_i[23] ) );
  AO22X1_RVT U4771 ( .A1(\read_value_mux[30][24] ), .A2(n3067), .A3(
        write_data[24]), .A4(n3066), .Y(\words[30]/data_i[24] ) );
  AO22X1_RVT U4772 ( .A1(\read_value_mux[30][25] ), .A2(n3067), .A3(
        write_data[25]), .A4(n3066), .Y(\words[30]/data_i[25] ) );
  AO22X1_RVT U4773 ( .A1(\read_value_mux[30][26] ), .A2(n3067), .A3(
        write_data[26]), .A4(n3066), .Y(\words[30]/data_i[26] ) );
  AO22X1_RVT U4774 ( .A1(\read_value_mux[30][27] ), .A2(n3067), .A3(
        write_data[27]), .A4(n3066), .Y(\words[30]/data_i[27] ) );
  AO22X1_RVT U4775 ( .A1(\read_value_mux[30][28] ), .A2(n3067), .A3(
        write_data[28]), .A4(n3066), .Y(\words[30]/data_i[28] ) );
  AO22X1_RVT U4776 ( .A1(\read_value_mux[30][29] ), .A2(n3067), .A3(
        write_data[29]), .A4(n3066), .Y(\words[30]/data_i[29] ) );
  AO22X1_RVT U4777 ( .A1(\read_value_mux[30][2] ), .A2(n3067), .A3(
        write_data[2]), .A4(n3066), .Y(\words[30]/data_i[2] ) );
  AO22X1_RVT U4778 ( .A1(n3066), .A2(write_data[30]), .A3(
        \read_value_mux[30][30] ), .A4(n3067), .Y(\words[30]/data_i[30] ) );
  AO22X1_RVT U4779 ( .A1(\read_value_mux[30][31] ), .A2(n3067), .A3(
        write_data[31]), .A4(n3066), .Y(\words[30]/data_i[31] ) );
  AO22X1_RVT U4780 ( .A1(\read_value_mux[30][3] ), .A2(n3067), .A3(
        write_data[3]), .A4(n3066), .Y(\words[30]/data_i[3] ) );
  AO22X1_RVT U4781 ( .A1(\read_value_mux[30][4] ), .A2(n3067), .A3(
        write_data[4]), .A4(n3066), .Y(\words[30]/data_i[4] ) );
  AO22X1_RVT U4782 ( .A1(\read_value_mux[30][5] ), .A2(n3067), .A3(
        write_data[5]), .A4(n3066), .Y(\words[30]/data_i[5] ) );
  AO22X1_RVT U4783 ( .A1(\read_value_mux[30][6] ), .A2(n3067), .A3(
        write_data[6]), .A4(n3066), .Y(\words[30]/data_i[6] ) );
  AO22X1_RVT U4784 ( .A1(\read_value_mux[30][7] ), .A2(n3067), .A3(
        write_data[7]), .A4(n3066), .Y(\words[30]/data_i[7] ) );
  AO22X1_RVT U4785 ( .A1(\read_value_mux[30][8] ), .A2(n3067), .A3(
        write_data[8]), .A4(n3066), .Y(\words[30]/data_i[8] ) );
  AO22X1_RVT U4786 ( .A1(\read_value_mux[30][9] ), .A2(n3067), .A3(
        write_data[9]), .A4(n3066), .Y(\words[30]/data_i[9] ) );
  AO21X1_RVT U4787 ( .A1(\words[30]/valid_o ), .A2(n3067), .A3(n3066), .Y(
        \words[30]/valid_i ) );
  AO22X1_RVT U4788 ( .A1(\read_value_mux[31][0] ), .A2(n3072), .A3(
        write_data[0]), .A4(n3071), .Y(\words[31]/data_i[0] ) );
  AO22X1_RVT U4789 ( .A1(\read_value_mux[31][10] ), .A2(n3072), .A3(
        write_data[10]), .A4(n3071), .Y(\words[31]/data_i[10] ) );
  AO22X1_RVT U4790 ( .A1(\read_value_mux[31][11] ), .A2(n3072), .A3(
        write_data[11]), .A4(n3071), .Y(\words[31]/data_i[11] ) );
  AO22X1_RVT U4791 ( .A1(\read_value_mux[31][12] ), .A2(n3072), .A3(
        write_data[12]), .A4(n3071), .Y(\words[31]/data_i[12] ) );
  AO22X1_RVT U4792 ( .A1(\read_value_mux[31][13] ), .A2(n3072), .A3(
        write_data[13]), .A4(n3071), .Y(\words[31]/data_i[13] ) );
  AO22X1_RVT U4793 ( .A1(\read_value_mux[31][14] ), .A2(n3072), .A3(
        write_data[14]), .A4(n3071), .Y(\words[31]/data_i[14] ) );
  AO22X1_RVT U4794 ( .A1(\read_value_mux[31][15] ), .A2(n3072), .A3(
        write_data[15]), .A4(n3071), .Y(\words[31]/data_i[15] ) );
  AO22X1_RVT U4795 ( .A1(\read_value_mux[31][16] ), .A2(n3072), .A3(
        write_data[16]), .A4(n3071), .Y(\words[31]/data_i[16] ) );
  AO22X1_RVT U4796 ( .A1(\read_value_mux[31][17] ), .A2(n3072), .A3(
        write_data[17]), .A4(n3071), .Y(\words[31]/data_i[17] ) );
  AO22X1_RVT U4797 ( .A1(\read_value_mux[31][18] ), .A2(n3072), .A3(
        write_data[18]), .A4(n3071), .Y(\words[31]/data_i[18] ) );
  AO22X1_RVT U4798 ( .A1(\read_value_mux[31][19] ), .A2(n3072), .A3(
        write_data[19]), .A4(n3071), .Y(\words[31]/data_i[19] ) );
  AO22X1_RVT U4799 ( .A1(n3071), .A2(write_data[1]), .A3(
        \read_value_mux[31][1] ), .A4(n3072), .Y(\words[31]/data_i[1] ) );
  AO22X1_RVT U4800 ( .A1(\read_value_mux[31][20] ), .A2(n3072), .A3(
        write_data[20]), .A4(n3071), .Y(\words[31]/data_i[20] ) );
  AO22X1_RVT U4801 ( .A1(\read_value_mux[31][21] ), .A2(n3072), .A3(
        write_data[21]), .A4(n3071), .Y(\words[31]/data_i[21] ) );
  AO22X1_RVT U4802 ( .A1(\read_value_mux[31][22] ), .A2(n3072), .A3(
        write_data[22]), .A4(n3071), .Y(\words[31]/data_i[22] ) );
  AO22X1_RVT U4803 ( .A1(\read_value_mux[31][23] ), .A2(n3072), .A3(
        write_data[23]), .A4(n3071), .Y(\words[31]/data_i[23] ) );
  AO22X1_RVT U4804 ( .A1(\read_value_mux[31][24] ), .A2(n3072), .A3(
        write_data[24]), .A4(n3071), .Y(\words[31]/data_i[24] ) );
  AO22X1_RVT U4805 ( .A1(\read_value_mux[31][25] ), .A2(n3072), .A3(
        write_data[25]), .A4(n3071), .Y(\words[31]/data_i[25] ) );
  AO22X1_RVT U4806 ( .A1(\read_value_mux[31][26] ), .A2(n3072), .A3(
        write_data[26]), .A4(n3071), .Y(\words[31]/data_i[26] ) );
  AO22X1_RVT U4807 ( .A1(\read_value_mux[31][27] ), .A2(n3072), .A3(
        write_data[27]), .A4(n3071), .Y(\words[31]/data_i[27] ) );
  AO22X1_RVT U4808 ( .A1(\read_value_mux[31][28] ), .A2(n3072), .A3(
        write_data[28]), .A4(n3071), .Y(\words[31]/data_i[28] ) );
  AO22X1_RVT U4809 ( .A1(\read_value_mux[31][29] ), .A2(n3072), .A3(
        write_data[29]), .A4(n3071), .Y(\words[31]/data_i[29] ) );
  AO22X1_RVT U4810 ( .A1(\read_value_mux[31][2] ), .A2(n3072), .A3(
        write_data[2]), .A4(n3071), .Y(\words[31]/data_i[2] ) );
  AO22X1_RVT U4811 ( .A1(n3071), .A2(write_data[30]), .A3(
        \read_value_mux[31][30] ), .A4(n3072), .Y(\words[31]/data_i[30] ) );
  AO22X1_RVT U4812 ( .A1(\read_value_mux[31][31] ), .A2(n3072), .A3(
        write_data[31]), .A4(n3071), .Y(\words[31]/data_i[31] ) );
  AO22X1_RVT U4813 ( .A1(\read_value_mux[31][3] ), .A2(n3072), .A3(
        write_data[3]), .A4(n3071), .Y(\words[31]/data_i[3] ) );
  AO22X1_RVT U4814 ( .A1(\read_value_mux[31][4] ), .A2(n3072), .A3(
        write_data[4]), .A4(n3071), .Y(\words[31]/data_i[4] ) );
  AO22X1_RVT U4815 ( .A1(\read_value_mux[31][5] ), .A2(n3072), .A3(
        write_data[5]), .A4(n3071), .Y(\words[31]/data_i[5] ) );
  AO22X1_RVT U4816 ( .A1(\read_value_mux[31][6] ), .A2(n3072), .A3(
        write_data[6]), .A4(n3071), .Y(\words[31]/data_i[6] ) );
  AO22X1_RVT U4817 ( .A1(\read_value_mux[31][7] ), .A2(n3072), .A3(
        write_data[7]), .A4(n3071), .Y(\words[31]/data_i[7] ) );
  AO22X1_RVT U4818 ( .A1(\read_value_mux[31][8] ), .A2(n3072), .A3(
        write_data[8]), .A4(n3071), .Y(\words[31]/data_i[8] ) );
  AO22X1_RVT U4819 ( .A1(\read_value_mux[31][9] ), .A2(n3072), .A3(
        write_data[9]), .A4(n3071), .Y(\words[31]/data_i[9] ) );
  AO21X1_RVT U4820 ( .A1(\words[31]/valid_o ), .A2(n3072), .A3(n3071), .Y(
        \words[31]/valid_i ) );
  AO22X1_RVT U4821 ( .A1(\read_value_mux[3][0] ), .A2(n3076), .A3(
        write_data[0]), .A4(n3075), .Y(\words[3]/data_i[0] ) );
  AO22X1_RVT U4822 ( .A1(\read_value_mux[3][10] ), .A2(n3076), .A3(
        write_data[10]), .A4(n3075), .Y(\words[3]/data_i[10] ) );
  AO22X1_RVT U4823 ( .A1(\read_value_mux[3][11] ), .A2(n3076), .A3(
        write_data[11]), .A4(n3075), .Y(\words[3]/data_i[11] ) );
  AO22X1_RVT U4824 ( .A1(\read_value_mux[3][12] ), .A2(n3076), .A3(
        write_data[12]), .A4(n3075), .Y(\words[3]/data_i[12] ) );
  AO22X1_RVT U4825 ( .A1(\read_value_mux[3][13] ), .A2(n3076), .A3(
        write_data[13]), .A4(n3075), .Y(\words[3]/data_i[13] ) );
  AO22X1_RVT U4826 ( .A1(\read_value_mux[3][14] ), .A2(n3076), .A3(
        write_data[14]), .A4(n3075), .Y(\words[3]/data_i[14] ) );
  AO22X1_RVT U4827 ( .A1(\read_value_mux[3][15] ), .A2(n3076), .A3(
        write_data[15]), .A4(n3075), .Y(\words[3]/data_i[15] ) );
  AO22X1_RVT U4828 ( .A1(\read_value_mux[3][16] ), .A2(n3076), .A3(
        write_data[16]), .A4(n3075), .Y(\words[3]/data_i[16] ) );
  AO22X1_RVT U4829 ( .A1(\read_value_mux[3][17] ), .A2(n3076), .A3(
        write_data[17]), .A4(n3075), .Y(\words[3]/data_i[17] ) );
  AO22X1_RVT U4830 ( .A1(\read_value_mux[3][18] ), .A2(n3076), .A3(
        write_data[18]), .A4(n3075), .Y(\words[3]/data_i[18] ) );
  AO22X1_RVT U4831 ( .A1(\read_value_mux[3][19] ), .A2(n3076), .A3(
        write_data[19]), .A4(n3075), .Y(\words[3]/data_i[19] ) );
  AO22X1_RVT U4832 ( .A1(n3075), .A2(write_data[1]), .A3(
        \read_value_mux[3][1] ), .A4(n3076), .Y(\words[3]/data_i[1] ) );
  AO22X1_RVT U4833 ( .A1(\read_value_mux[3][20] ), .A2(n3076), .A3(
        write_data[20]), .A4(n3075), .Y(\words[3]/data_i[20] ) );
  AO22X1_RVT U4834 ( .A1(\read_value_mux[3][21] ), .A2(n3076), .A3(
        write_data[21]), .A4(n3075), .Y(\words[3]/data_i[21] ) );
  AO22X1_RVT U4835 ( .A1(\read_value_mux[3][22] ), .A2(n3076), .A3(
        write_data[22]), .A4(n3075), .Y(\words[3]/data_i[22] ) );
  AO22X1_RVT U4836 ( .A1(\read_value_mux[3][23] ), .A2(n3076), .A3(
        write_data[23]), .A4(n3075), .Y(\words[3]/data_i[23] ) );
  AO22X1_RVT U4837 ( .A1(\read_value_mux[3][24] ), .A2(n3076), .A3(
        write_data[24]), .A4(n3075), .Y(\words[3]/data_i[24] ) );
  AO22X1_RVT U4838 ( .A1(\read_value_mux[3][25] ), .A2(n3076), .A3(
        write_data[25]), .A4(n3075), .Y(\words[3]/data_i[25] ) );
  AO22X1_RVT U4839 ( .A1(\read_value_mux[3][26] ), .A2(n3076), .A3(
        write_data[26]), .A4(n3075), .Y(\words[3]/data_i[26] ) );
  AO22X1_RVT U4840 ( .A1(\read_value_mux[3][27] ), .A2(n3076), .A3(
        write_data[27]), .A4(n3075), .Y(\words[3]/data_i[27] ) );
  AO22X1_RVT U4841 ( .A1(\read_value_mux[3][28] ), .A2(n3076), .A3(
        write_data[28]), .A4(n3075), .Y(\words[3]/data_i[28] ) );
  AO22X1_RVT U4842 ( .A1(\read_value_mux[3][29] ), .A2(n3076), .A3(
        write_data[29]), .A4(n3075), .Y(\words[3]/data_i[29] ) );
  AO22X1_RVT U4843 ( .A1(\read_value_mux[3][2] ), .A2(n3076), .A3(
        write_data[2]), .A4(n3075), .Y(\words[3]/data_i[2] ) );
  AO22X1_RVT U4844 ( .A1(n3075), .A2(write_data[30]), .A3(
        \read_value_mux[3][30] ), .A4(n3076), .Y(\words[3]/data_i[30] ) );
  AO22X1_RVT U4845 ( .A1(\read_value_mux[3][31] ), .A2(n3076), .A3(
        write_data[31]), .A4(n3075), .Y(\words[3]/data_i[31] ) );
  AO22X1_RVT U4846 ( .A1(\read_value_mux[3][3] ), .A2(n3076), .A3(
        write_data[3]), .A4(n3075), .Y(\words[3]/data_i[3] ) );
  AO22X1_RVT U4847 ( .A1(\read_value_mux[3][4] ), .A2(n3076), .A3(
        write_data[4]), .A4(n3075), .Y(\words[3]/data_i[4] ) );
  AO22X1_RVT U4848 ( .A1(\read_value_mux[3][5] ), .A2(n3076), .A3(
        write_data[5]), .A4(n3075), .Y(\words[3]/data_i[5] ) );
  AO22X1_RVT U4849 ( .A1(\read_value_mux[3][6] ), .A2(n3076), .A3(
        write_data[6]), .A4(n3075), .Y(\words[3]/data_i[6] ) );
  AO22X1_RVT U4850 ( .A1(\read_value_mux[3][7] ), .A2(n3076), .A3(
        write_data[7]), .A4(n3075), .Y(\words[3]/data_i[7] ) );
  AO22X1_RVT U4851 ( .A1(\read_value_mux[3][8] ), .A2(n3076), .A3(
        write_data[8]), .A4(n3075), .Y(\words[3]/data_i[8] ) );
  AO22X1_RVT U4852 ( .A1(\read_value_mux[3][9] ), .A2(n3076), .A3(
        write_data[9]), .A4(n3075), .Y(\words[3]/data_i[9] ) );
  AO21X1_RVT U4853 ( .A1(\words[3]/valid_o ), .A2(n3076), .A3(n3075), .Y(
        \words[3]/valid_i ) );
  AO22X1_RVT U4854 ( .A1(\read_value_mux[4][0] ), .A2(n1679), .A3(
        write_data[0]), .A4(n3077), .Y(\words[4]/data_i[0] ) );
  AO22X1_RVT U4855 ( .A1(\read_value_mux[4][10] ), .A2(n1679), .A3(
        write_data[10]), .A4(n3077), .Y(\words[4]/data_i[10] ) );
  AO22X1_RVT U4856 ( .A1(\read_value_mux[4][11] ), .A2(n1679), .A3(
        write_data[11]), .A4(n3077), .Y(\words[4]/data_i[11] ) );
  AO22X1_RVT U4857 ( .A1(\read_value_mux[4][12] ), .A2(n1679), .A3(
        write_data[12]), .A4(n3077), .Y(\words[4]/data_i[12] ) );
  AO22X1_RVT U4858 ( .A1(\read_value_mux[4][13] ), .A2(n1679), .A3(
        write_data[13]), .A4(n3077), .Y(\words[4]/data_i[13] ) );
  AO22X1_RVT U4859 ( .A1(\read_value_mux[4][14] ), .A2(n1679), .A3(
        write_data[14]), .A4(n3077), .Y(\words[4]/data_i[14] ) );
  AO22X1_RVT U4860 ( .A1(\read_value_mux[4][15] ), .A2(n1679), .A3(
        write_data[15]), .A4(n3077), .Y(\words[4]/data_i[15] ) );
  AO22X1_RVT U4861 ( .A1(\read_value_mux[4][16] ), .A2(n1679), .A3(
        write_data[16]), .A4(n3077), .Y(\words[4]/data_i[16] ) );
  AO22X1_RVT U4862 ( .A1(\read_value_mux[4][17] ), .A2(n1679), .A3(
        write_data[17]), .A4(n3077), .Y(\words[4]/data_i[17] ) );
  AO22X1_RVT U4863 ( .A1(\read_value_mux[4][18] ), .A2(n1679), .A3(
        write_data[18]), .A4(n3077), .Y(\words[4]/data_i[18] ) );
  AO22X1_RVT U4864 ( .A1(\read_value_mux[4][19] ), .A2(n1679), .A3(
        write_data[19]), .A4(n3077), .Y(\words[4]/data_i[19] ) );
  AO22X1_RVT U4865 ( .A1(n3077), .A2(write_data[1]), .A3(
        \read_value_mux[4][1] ), .A4(n1679), .Y(\words[4]/data_i[1] ) );
  AO22X1_RVT U4866 ( .A1(\read_value_mux[4][20] ), .A2(n1679), .A3(
        write_data[20]), .A4(n3077), .Y(\words[4]/data_i[20] ) );
  AO22X1_RVT U4867 ( .A1(\read_value_mux[4][21] ), .A2(n1679), .A3(
        write_data[21]), .A4(n3077), .Y(\words[4]/data_i[21] ) );
  AO22X1_RVT U4868 ( .A1(\read_value_mux[4][22] ), .A2(n1679), .A3(
        write_data[22]), .A4(n3077), .Y(\words[4]/data_i[22] ) );
  AO22X1_RVT U4869 ( .A1(\read_value_mux[4][23] ), .A2(n1679), .A3(
        write_data[23]), .A4(n3077), .Y(\words[4]/data_i[23] ) );
  AO22X1_RVT U4870 ( .A1(\read_value_mux[4][24] ), .A2(n1679), .A3(
        write_data[24]), .A4(n3077), .Y(\words[4]/data_i[24] ) );
  AO22X1_RVT U4871 ( .A1(\read_value_mux[4][25] ), .A2(n1679), .A3(
        write_data[25]), .A4(n3077), .Y(\words[4]/data_i[25] ) );
  AO22X1_RVT U4872 ( .A1(\read_value_mux[4][26] ), .A2(n1679), .A3(
        write_data[26]), .A4(n3077), .Y(\words[4]/data_i[26] ) );
  AO22X1_RVT U4873 ( .A1(\read_value_mux[4][27] ), .A2(n1679), .A3(
        write_data[27]), .A4(n3077), .Y(\words[4]/data_i[27] ) );
  AO22X1_RVT U4874 ( .A1(\read_value_mux[4][28] ), .A2(n1679), .A3(
        write_data[28]), .A4(n3077), .Y(\words[4]/data_i[28] ) );
  AO22X1_RVT U4875 ( .A1(\read_value_mux[4][29] ), .A2(n1679), .A3(
        write_data[29]), .A4(n3077), .Y(\words[4]/data_i[29] ) );
  AO22X1_RVT U4876 ( .A1(\read_value_mux[4][2] ), .A2(n1679), .A3(
        write_data[2]), .A4(n3077), .Y(\words[4]/data_i[2] ) );
  AO22X1_RVT U4877 ( .A1(n3077), .A2(write_data[30]), .A3(
        \read_value_mux[4][30] ), .A4(n1679), .Y(\words[4]/data_i[30] ) );
  AO22X1_RVT U4878 ( .A1(\read_value_mux[4][31] ), .A2(n1679), .A3(
        write_data[31]), .A4(n3077), .Y(\words[4]/data_i[31] ) );
  AO22X1_RVT U4879 ( .A1(\read_value_mux[4][3] ), .A2(n1679), .A3(
        write_data[3]), .A4(n3077), .Y(\words[4]/data_i[3] ) );
  AO22X1_RVT U4880 ( .A1(\read_value_mux[4][4] ), .A2(n1679), .A3(
        write_data[4]), .A4(n3077), .Y(\words[4]/data_i[4] ) );
  AO22X1_RVT U4881 ( .A1(\read_value_mux[4][5] ), .A2(n1679), .A3(
        write_data[5]), .A4(n3077), .Y(\words[4]/data_i[5] ) );
  AO22X1_RVT U4882 ( .A1(\read_value_mux[4][6] ), .A2(n1679), .A3(
        write_data[6]), .A4(n3077), .Y(\words[4]/data_i[6] ) );
  AO22X1_RVT U4883 ( .A1(\read_value_mux[4][7] ), .A2(n1679), .A3(
        write_data[7]), .A4(n3077), .Y(\words[4]/data_i[7] ) );
  AO22X1_RVT U4884 ( .A1(\read_value_mux[4][8] ), .A2(n1679), .A3(
        write_data[8]), .A4(n3077), .Y(\words[4]/data_i[8] ) );
  AO22X1_RVT U4885 ( .A1(\read_value_mux[4][9] ), .A2(n1679), .A3(
        write_data[9]), .A4(n3077), .Y(\words[4]/data_i[9] ) );
  AO21X1_RVT U4886 ( .A1(\words[4]/valid_o ), .A2(n1679), .A3(n3077), .Y(
        \words[4]/valid_i ) );
  AO22X1_RVT U4887 ( .A1(\read_value_mux[5][0] ), .A2(n1684), .A3(
        write_data[0]), .A4(n3078), .Y(\words[5]/data_i[0] ) );
  AO22X1_RVT U4888 ( .A1(\read_value_mux[5][10] ), .A2(n1684), .A3(
        write_data[10]), .A4(n3078), .Y(\words[5]/data_i[10] ) );
  AO22X1_RVT U4889 ( .A1(\read_value_mux[5][11] ), .A2(n1684), .A3(
        write_data[11]), .A4(n3078), .Y(\words[5]/data_i[11] ) );
  AO22X1_RVT U4890 ( .A1(\read_value_mux[5][12] ), .A2(n1684), .A3(
        write_data[12]), .A4(n3078), .Y(\words[5]/data_i[12] ) );
  AO22X1_RVT U4891 ( .A1(\read_value_mux[5][13] ), .A2(n1684), .A3(
        write_data[13]), .A4(n3078), .Y(\words[5]/data_i[13] ) );
  AO22X1_RVT U4892 ( .A1(\read_value_mux[5][14] ), .A2(n1684), .A3(
        write_data[14]), .A4(n3078), .Y(\words[5]/data_i[14] ) );
  AO22X1_RVT U4893 ( .A1(\read_value_mux[5][15] ), .A2(n1684), .A3(
        write_data[15]), .A4(n3078), .Y(\words[5]/data_i[15] ) );
  AO22X1_RVT U4894 ( .A1(\read_value_mux[5][16] ), .A2(n1684), .A3(
        write_data[16]), .A4(n3078), .Y(\words[5]/data_i[16] ) );
  AO22X1_RVT U4895 ( .A1(\read_value_mux[5][17] ), .A2(n1684), .A3(
        write_data[17]), .A4(n3078), .Y(\words[5]/data_i[17] ) );
  AO22X1_RVT U4896 ( .A1(\read_value_mux[5][18] ), .A2(n1684), .A3(
        write_data[18]), .A4(n3078), .Y(\words[5]/data_i[18] ) );
  AO22X1_RVT U4897 ( .A1(\read_value_mux[5][19] ), .A2(n1684), .A3(
        write_data[19]), .A4(n3078), .Y(\words[5]/data_i[19] ) );
  AO22X1_RVT U4898 ( .A1(n3078), .A2(write_data[1]), .A3(
        \read_value_mux[5][1] ), .A4(n1684), .Y(\words[5]/data_i[1] ) );
  AO22X1_RVT U4899 ( .A1(\read_value_mux[5][20] ), .A2(n1684), .A3(
        write_data[20]), .A4(n3078), .Y(\words[5]/data_i[20] ) );
  AO22X1_RVT U4900 ( .A1(\read_value_mux[5][21] ), .A2(n1684), .A3(
        write_data[21]), .A4(n3078), .Y(\words[5]/data_i[21] ) );
  AO22X1_RVT U4901 ( .A1(\read_value_mux[5][22] ), .A2(n1684), .A3(
        write_data[22]), .A4(n3078), .Y(\words[5]/data_i[22] ) );
  AO22X1_RVT U4902 ( .A1(\read_value_mux[5][23] ), .A2(n1684), .A3(
        write_data[23]), .A4(n3078), .Y(\words[5]/data_i[23] ) );
  AO22X1_RVT U4903 ( .A1(\read_value_mux[5][24] ), .A2(n1684), .A3(
        write_data[24]), .A4(n3078), .Y(\words[5]/data_i[24] ) );
  AO22X1_RVT U4904 ( .A1(\read_value_mux[5][25] ), .A2(n1684), .A3(
        write_data[25]), .A4(n3078), .Y(\words[5]/data_i[25] ) );
  AO22X1_RVT U4905 ( .A1(\read_value_mux[5][26] ), .A2(n1684), .A3(
        write_data[26]), .A4(n3078), .Y(\words[5]/data_i[26] ) );
  AO22X1_RVT U4906 ( .A1(\read_value_mux[5][27] ), .A2(n1684), .A3(
        write_data[27]), .A4(n3078), .Y(\words[5]/data_i[27] ) );
  AO22X1_RVT U4907 ( .A1(\read_value_mux[5][28] ), .A2(n1684), .A3(
        write_data[28]), .A4(n3078), .Y(\words[5]/data_i[28] ) );
  AO22X1_RVT U4908 ( .A1(\read_value_mux[5][29] ), .A2(n1684), .A3(
        write_data[29]), .A4(n3078), .Y(\words[5]/data_i[29] ) );
  AO22X1_RVT U4909 ( .A1(\read_value_mux[5][2] ), .A2(n1684), .A3(
        write_data[2]), .A4(n3078), .Y(\words[5]/data_i[2] ) );
  AO22X1_RVT U4910 ( .A1(n3078), .A2(write_data[30]), .A3(
        \read_value_mux[5][30] ), .A4(n1684), .Y(\words[5]/data_i[30] ) );
  AO22X1_RVT U4911 ( .A1(\read_value_mux[5][31] ), .A2(n1684), .A3(
        write_data[31]), .A4(n3078), .Y(\words[5]/data_i[31] ) );
  AO22X1_RVT U4912 ( .A1(\read_value_mux[5][3] ), .A2(n1684), .A3(
        write_data[3]), .A4(n3078), .Y(\words[5]/data_i[3] ) );
  AO22X1_RVT U4913 ( .A1(\read_value_mux[5][4] ), .A2(n1684), .A3(
        write_data[4]), .A4(n3078), .Y(\words[5]/data_i[4] ) );
  AO22X1_RVT U4914 ( .A1(\read_value_mux[5][5] ), .A2(n1684), .A3(
        write_data[5]), .A4(n3078), .Y(\words[5]/data_i[5] ) );
  AO22X1_RVT U4915 ( .A1(\read_value_mux[5][6] ), .A2(n1684), .A3(
        write_data[6]), .A4(n3078), .Y(\words[5]/data_i[6] ) );
  AO22X1_RVT U4916 ( .A1(\read_value_mux[5][7] ), .A2(n1684), .A3(
        write_data[7]), .A4(n3078), .Y(\words[5]/data_i[7] ) );
  AO22X1_RVT U4917 ( .A1(\read_value_mux[5][8] ), .A2(n1684), .A3(
        write_data[8]), .A4(n3078), .Y(\words[5]/data_i[8] ) );
  AO22X1_RVT U4918 ( .A1(\read_value_mux[5][9] ), .A2(n1684), .A3(
        write_data[9]), .A4(n3078), .Y(\words[5]/data_i[9] ) );
  AO21X1_RVT U4919 ( .A1(\words[5]/valid_o ), .A2(n1684), .A3(n3078), .Y(
        \words[5]/valid_i ) );
  AO22X1_RVT U4920 ( .A1(\read_value_mux[6][0] ), .A2(n3082), .A3(
        write_data[0]), .A4(n3081), .Y(\words[6]/data_i[0] ) );
  AO22X1_RVT U4921 ( .A1(\read_value_mux[6][10] ), .A2(n3082), .A3(
        write_data[10]), .A4(n3081), .Y(\words[6]/data_i[10] ) );
  AO22X1_RVT U4922 ( .A1(\read_value_mux[6][11] ), .A2(n3082), .A3(
        write_data[11]), .A4(n3081), .Y(\words[6]/data_i[11] ) );
  AO22X1_RVT U4923 ( .A1(\read_value_mux[6][12] ), .A2(n3082), .A3(
        write_data[12]), .A4(n3081), .Y(\words[6]/data_i[12] ) );
  AO22X1_RVT U4924 ( .A1(\read_value_mux[6][13] ), .A2(n3082), .A3(
        write_data[13]), .A4(n3081), .Y(\words[6]/data_i[13] ) );
  AO22X1_RVT U4925 ( .A1(\read_value_mux[6][14] ), .A2(n3082), .A3(
        write_data[14]), .A4(n3081), .Y(\words[6]/data_i[14] ) );
  AO22X1_RVT U4926 ( .A1(\read_value_mux[6][15] ), .A2(n3082), .A3(
        write_data[15]), .A4(n3081), .Y(\words[6]/data_i[15] ) );
  AO22X1_RVT U4927 ( .A1(\read_value_mux[6][16] ), .A2(n3082), .A3(
        write_data[16]), .A4(n3081), .Y(\words[6]/data_i[16] ) );
  AO22X1_RVT U4928 ( .A1(\read_value_mux[6][17] ), .A2(n3082), .A3(
        write_data[17]), .A4(n3081), .Y(\words[6]/data_i[17] ) );
  AO22X1_RVT U4929 ( .A1(\read_value_mux[6][18] ), .A2(n3082), .A3(
        write_data[18]), .A4(n3081), .Y(\words[6]/data_i[18] ) );
  AO22X1_RVT U4930 ( .A1(\read_value_mux[6][19] ), .A2(n3082), .A3(
        write_data[19]), .A4(n3081), .Y(\words[6]/data_i[19] ) );
  AO22X1_RVT U4931 ( .A1(n3081), .A2(write_data[1]), .A3(
        \read_value_mux[6][1] ), .A4(n3082), .Y(\words[6]/data_i[1] ) );
  AO22X1_RVT U4932 ( .A1(\read_value_mux[6][20] ), .A2(n3082), .A3(
        write_data[20]), .A4(n3081), .Y(\words[6]/data_i[20] ) );
  AO22X1_RVT U4933 ( .A1(\read_value_mux[6][21] ), .A2(n3082), .A3(
        write_data[21]), .A4(n3081), .Y(\words[6]/data_i[21] ) );
  AO22X1_RVT U4934 ( .A1(\read_value_mux[6][22] ), .A2(n3082), .A3(
        write_data[22]), .A4(n3081), .Y(\words[6]/data_i[22] ) );
  AO22X1_RVT U4935 ( .A1(\read_value_mux[6][23] ), .A2(n3082), .A3(
        write_data[23]), .A4(n3081), .Y(\words[6]/data_i[23] ) );
  AO22X1_RVT U4936 ( .A1(\read_value_mux[6][24] ), .A2(n3082), .A3(
        write_data[24]), .A4(n3081), .Y(\words[6]/data_i[24] ) );
  AO22X1_RVT U4937 ( .A1(\read_value_mux[6][25] ), .A2(n3082), .A3(
        write_data[25]), .A4(n3081), .Y(\words[6]/data_i[25] ) );
  AO22X1_RVT U4938 ( .A1(\read_value_mux[6][26] ), .A2(n3082), .A3(
        write_data[26]), .A4(n3081), .Y(\words[6]/data_i[26] ) );
  AO22X1_RVT U4939 ( .A1(\read_value_mux[6][27] ), .A2(n3082), .A3(
        write_data[27]), .A4(n3081), .Y(\words[6]/data_i[27] ) );
  AO22X1_RVT U4940 ( .A1(\read_value_mux[6][28] ), .A2(n3082), .A3(
        write_data[28]), .A4(n3081), .Y(\words[6]/data_i[28] ) );
  AO22X1_RVT U4941 ( .A1(\read_value_mux[6][29] ), .A2(n3082), .A3(
        write_data[29]), .A4(n3081), .Y(\words[6]/data_i[29] ) );
  AO22X1_RVT U4942 ( .A1(\read_value_mux[6][2] ), .A2(n3082), .A3(
        write_data[2]), .A4(n3081), .Y(\words[6]/data_i[2] ) );
  AO22X1_RVT U4943 ( .A1(n3081), .A2(write_data[30]), .A3(
        \read_value_mux[6][30] ), .A4(n3082), .Y(\words[6]/data_i[30] ) );
  AO22X1_RVT U4944 ( .A1(\read_value_mux[6][31] ), .A2(n3082), .A3(
        write_data[31]), .A4(n3081), .Y(\words[6]/data_i[31] ) );
  AO22X1_RVT U4945 ( .A1(\read_value_mux[6][3] ), .A2(n3082), .A3(
        write_data[3]), .A4(n3081), .Y(\words[6]/data_i[3] ) );
  AO22X1_RVT U4946 ( .A1(\read_value_mux[6][4] ), .A2(n3082), .A3(
        write_data[4]), .A4(n3081), .Y(\words[6]/data_i[4] ) );
  AO22X1_RVT U4947 ( .A1(\read_value_mux[6][5] ), .A2(n3082), .A3(
        write_data[5]), .A4(n3081), .Y(\words[6]/data_i[5] ) );
  AO22X1_RVT U4948 ( .A1(\read_value_mux[6][6] ), .A2(n3082), .A3(
        write_data[6]), .A4(n3081), .Y(\words[6]/data_i[6] ) );
  AO22X1_RVT U4949 ( .A1(\read_value_mux[6][7] ), .A2(n3082), .A3(
        write_data[7]), .A4(n3081), .Y(\words[6]/data_i[7] ) );
  AO22X1_RVT U4950 ( .A1(\read_value_mux[6][8] ), .A2(n3082), .A3(
        write_data[8]), .A4(n3081), .Y(\words[6]/data_i[8] ) );
  AO22X1_RVT U4951 ( .A1(\read_value_mux[6][9] ), .A2(n3082), .A3(
        write_data[9]), .A4(n3081), .Y(\words[6]/data_i[9] ) );
  AO21X1_RVT U4952 ( .A1(\words[6]/valid_o ), .A2(n3082), .A3(n3081), .Y(
        \words[6]/valid_i ) );
  AO22X1_RVT U4953 ( .A1(\read_value_mux[7][0] ), .A2(n1634), .A3(
        write_data[0]), .A4(n3089), .Y(\words[7]/data_i[0] ) );
  AO22X1_RVT U4954 ( .A1(\read_value_mux[7][10] ), .A2(n1634), .A3(
        write_data[10]), .A4(n3089), .Y(\words[7]/data_i[10] ) );
  AO22X1_RVT U4955 ( .A1(\read_value_mux[7][11] ), .A2(n1634), .A3(
        write_data[11]), .A4(n3089), .Y(\words[7]/data_i[11] ) );
  AO22X1_RVT U4956 ( .A1(\read_value_mux[7][12] ), .A2(n1634), .A3(
        write_data[12]), .A4(n3089), .Y(\words[7]/data_i[12] ) );
  AO22X1_RVT U4957 ( .A1(\read_value_mux[7][13] ), .A2(n1634), .A3(
        write_data[13]), .A4(n3089), .Y(\words[7]/data_i[13] ) );
  AO22X1_RVT U4958 ( .A1(\read_value_mux[7][14] ), .A2(n1634), .A3(
        write_data[14]), .A4(n3089), .Y(\words[7]/data_i[14] ) );
  AO22X1_RVT U4959 ( .A1(\read_value_mux[7][15] ), .A2(n1634), .A3(
        write_data[15]), .A4(n3089), .Y(\words[7]/data_i[15] ) );
  AO22X1_RVT U4960 ( .A1(\read_value_mux[7][16] ), .A2(n1634), .A3(
        write_data[16]), .A4(n3089), .Y(\words[7]/data_i[16] ) );
  AO22X1_RVT U4961 ( .A1(\read_value_mux[7][17] ), .A2(n1634), .A3(
        write_data[17]), .A4(n3089), .Y(\words[7]/data_i[17] ) );
  AO22X1_RVT U4962 ( .A1(\read_value_mux[7][18] ), .A2(n1634), .A3(
        write_data[18]), .A4(n3089), .Y(\words[7]/data_i[18] ) );
  AO22X1_RVT U4963 ( .A1(\read_value_mux[7][19] ), .A2(n1634), .A3(
        write_data[19]), .A4(n3089), .Y(\words[7]/data_i[19] ) );
  AO22X1_RVT U4964 ( .A1(n3089), .A2(write_data[1]), .A3(
        \read_value_mux[7][1] ), .A4(n1634), .Y(\words[7]/data_i[1] ) );
  AO22X1_RVT U4965 ( .A1(\read_value_mux[7][20] ), .A2(n1634), .A3(
        write_data[20]), .A4(n3089), .Y(\words[7]/data_i[20] ) );
  AO22X1_RVT U4966 ( .A1(\read_value_mux[7][21] ), .A2(n1634), .A3(
        write_data[21]), .A4(n3089), .Y(\words[7]/data_i[21] ) );
  AO22X1_RVT U4967 ( .A1(\read_value_mux[7][22] ), .A2(n1634), .A3(
        write_data[22]), .A4(n3089), .Y(\words[7]/data_i[22] ) );
  AO22X1_RVT U4968 ( .A1(\read_value_mux[7][23] ), .A2(n1634), .A3(
        write_data[23]), .A4(n3089), .Y(\words[7]/data_i[23] ) );
  AO22X1_RVT U4969 ( .A1(\read_value_mux[7][24] ), .A2(n1634), .A3(
        write_data[24]), .A4(n3089), .Y(\words[7]/data_i[24] ) );
  AO22X1_RVT U4970 ( .A1(\read_value_mux[7][25] ), .A2(n1634), .A3(
        write_data[25]), .A4(n3089), .Y(\words[7]/data_i[25] ) );
  AO22X1_RVT U4971 ( .A1(\read_value_mux[7][26] ), .A2(n1634), .A3(
        write_data[26]), .A4(n3089), .Y(\words[7]/data_i[26] ) );
  AO22X1_RVT U4972 ( .A1(\read_value_mux[7][27] ), .A2(n1634), .A3(
        write_data[27]), .A4(n3089), .Y(\words[7]/data_i[27] ) );
  AO22X1_RVT U4973 ( .A1(\read_value_mux[7][28] ), .A2(n1634), .A3(
        write_data[28]), .A4(n3089), .Y(\words[7]/data_i[28] ) );
  AO22X1_RVT U4974 ( .A1(\read_value_mux[7][29] ), .A2(n1634), .A3(
        write_data[29]), .A4(n3089), .Y(\words[7]/data_i[29] ) );
  AO22X1_RVT U4975 ( .A1(\read_value_mux[7][2] ), .A2(n1634), .A3(
        write_data[2]), .A4(n3089), .Y(\words[7]/data_i[2] ) );
  AO22X1_RVT U4976 ( .A1(n3089), .A2(write_data[30]), .A3(
        \read_value_mux[7][30] ), .A4(n1634), .Y(\words[7]/data_i[30] ) );
  AO22X1_RVT U4977 ( .A1(\read_value_mux[7][31] ), .A2(n1634), .A3(
        write_data[31]), .A4(n3089), .Y(\words[7]/data_i[31] ) );
  AO22X1_RVT U4978 ( .A1(\read_value_mux[7][3] ), .A2(n1634), .A3(
        write_data[3]), .A4(n3089), .Y(\words[7]/data_i[3] ) );
  AO22X1_RVT U4979 ( .A1(\read_value_mux[7][4] ), .A2(n1634), .A3(
        write_data[4]), .A4(n3089), .Y(\words[7]/data_i[4] ) );
  AO22X1_RVT U4980 ( .A1(\read_value_mux[7][5] ), .A2(n1634), .A3(
        write_data[5]), .A4(n3089), .Y(\words[7]/data_i[5] ) );
  AO22X1_RVT U4981 ( .A1(\read_value_mux[7][6] ), .A2(n1634), .A3(
        write_data[6]), .A4(n3089), .Y(\words[7]/data_i[6] ) );
  AO22X1_RVT U4982 ( .A1(\read_value_mux[7][7] ), .A2(n1634), .A3(
        write_data[7]), .A4(n3089), .Y(\words[7]/data_i[7] ) );
  AO22X1_RVT U4983 ( .A1(\read_value_mux[7][8] ), .A2(n1634), .A3(
        write_data[8]), .A4(n3089), .Y(\words[7]/data_i[8] ) );
  AO22X1_RVT U4984 ( .A1(\read_value_mux[7][9] ), .A2(n1634), .A3(
        write_data[9]), .A4(n3089), .Y(\words[7]/data_i[9] ) );
  AO21X1_RVT U4985 ( .A1(\words[7]/valid_o ), .A2(n1634), .A3(n3089), .Y(
        \words[7]/valid_i ) );
  AO22X1_RVT U4986 ( .A1(\read_value_mux[8][0] ), .A2(n1680), .A3(
        write_data[0]), .A4(n3092), .Y(\words[8]/data_i[0] ) );
  AO22X1_RVT U4987 ( .A1(\read_value_mux[8][10] ), .A2(n1680), .A3(
        write_data[10]), .A4(n3092), .Y(\words[8]/data_i[10] ) );
  AO22X1_RVT U4988 ( .A1(\read_value_mux[8][11] ), .A2(n1680), .A3(
        write_data[11]), .A4(n3092), .Y(\words[8]/data_i[11] ) );
  AO22X1_RVT U4989 ( .A1(\read_value_mux[8][12] ), .A2(n1680), .A3(
        write_data[12]), .A4(n3092), .Y(\words[8]/data_i[12] ) );
  AO22X1_RVT U4990 ( .A1(\read_value_mux[8][13] ), .A2(n1680), .A3(
        write_data[13]), .A4(n3092), .Y(\words[8]/data_i[13] ) );
  AO22X1_RVT U4991 ( .A1(\read_value_mux[8][14] ), .A2(n1680), .A3(
        write_data[14]), .A4(n3092), .Y(\words[8]/data_i[14] ) );
  AO22X1_RVT U4992 ( .A1(\read_value_mux[8][15] ), .A2(n1680), .A3(
        write_data[15]), .A4(n3092), .Y(\words[8]/data_i[15] ) );
  AO22X1_RVT U4993 ( .A1(\read_value_mux[8][16] ), .A2(n1680), .A3(
        write_data[16]), .A4(n3092), .Y(\words[8]/data_i[16] ) );
  AO22X1_RVT U4994 ( .A1(\read_value_mux[8][17] ), .A2(n1680), .A3(
        write_data[17]), .A4(n3092), .Y(\words[8]/data_i[17] ) );
  AO22X1_RVT U4995 ( .A1(\read_value_mux[8][18] ), .A2(n1680), .A3(
        write_data[18]), .A4(n3092), .Y(\words[8]/data_i[18] ) );
  AO22X1_RVT U4996 ( .A1(\read_value_mux[8][19] ), .A2(n1680), .A3(
        write_data[19]), .A4(n3092), .Y(\words[8]/data_i[19] ) );
  AO22X1_RVT U4997 ( .A1(n3092), .A2(write_data[1]), .A3(
        \read_value_mux[8][1] ), .A4(n1680), .Y(\words[8]/data_i[1] ) );
  AO22X1_RVT U4998 ( .A1(\read_value_mux[8][20] ), .A2(n1680), .A3(
        write_data[20]), .A4(n3092), .Y(\words[8]/data_i[20] ) );
  AO22X1_RVT U4999 ( .A1(\read_value_mux[8][21] ), .A2(n1680), .A3(
        write_data[21]), .A4(n3092), .Y(\words[8]/data_i[21] ) );
  AO22X1_RVT U5000 ( .A1(\read_value_mux[8][22] ), .A2(n1680), .A3(
        write_data[22]), .A4(n3092), .Y(\words[8]/data_i[22] ) );
  AO22X1_RVT U5001 ( .A1(\read_value_mux[8][23] ), .A2(n1680), .A3(
        write_data[23]), .A4(n3092), .Y(\words[8]/data_i[23] ) );
  AO22X1_RVT U5002 ( .A1(\read_value_mux[8][24] ), .A2(n1680), .A3(
        write_data[24]), .A4(n3092), .Y(\words[8]/data_i[24] ) );
  AO22X1_RVT U5003 ( .A1(\read_value_mux[8][25] ), .A2(n1680), .A3(
        write_data[25]), .A4(n3092), .Y(\words[8]/data_i[25] ) );
  AO22X1_RVT U5004 ( .A1(\read_value_mux[8][26] ), .A2(n1680), .A3(
        write_data[26]), .A4(n3092), .Y(\words[8]/data_i[26] ) );
  AO22X1_RVT U5005 ( .A1(\read_value_mux[8][27] ), .A2(n1680), .A3(
        write_data[27]), .A4(n3092), .Y(\words[8]/data_i[27] ) );
  AO22X1_RVT U5006 ( .A1(\read_value_mux[8][28] ), .A2(n1680), .A3(
        write_data[28]), .A4(n3092), .Y(\words[8]/data_i[28] ) );
  AO22X1_RVT U5007 ( .A1(\read_value_mux[8][29] ), .A2(n1680), .A3(
        write_data[29]), .A4(n3092), .Y(\words[8]/data_i[29] ) );
  AO22X1_RVT U5008 ( .A1(\read_value_mux[8][2] ), .A2(n1680), .A3(
        write_data[2]), .A4(n3092), .Y(\words[8]/data_i[2] ) );
  AO22X1_RVT U5009 ( .A1(n3092), .A2(write_data[30]), .A3(
        \read_value_mux[8][30] ), .A4(n1680), .Y(\words[8]/data_i[30] ) );
  AO22X1_RVT U5010 ( .A1(\read_value_mux[8][31] ), .A2(n1680), .A3(
        write_data[31]), .A4(n3092), .Y(\words[8]/data_i[31] ) );
  AO22X1_RVT U5011 ( .A1(\read_value_mux[8][3] ), .A2(n1680), .A3(
        write_data[3]), .A4(n3092), .Y(\words[8]/data_i[3] ) );
  AO22X1_RVT U5012 ( .A1(\read_value_mux[8][4] ), .A2(n1680), .A3(
        write_data[4]), .A4(n3092), .Y(\words[8]/data_i[4] ) );
  AO22X1_RVT U5013 ( .A1(\read_value_mux[8][5] ), .A2(n1680), .A3(
        write_data[5]), .A4(n3092), .Y(\words[8]/data_i[5] ) );
  AO22X1_RVT U5014 ( .A1(\read_value_mux[8][6] ), .A2(n1680), .A3(
        write_data[6]), .A4(n3092), .Y(\words[8]/data_i[6] ) );
  AO22X1_RVT U5015 ( .A1(\read_value_mux[8][7] ), .A2(n1680), .A3(
        write_data[7]), .A4(n3092), .Y(\words[8]/data_i[7] ) );
  AO22X1_RVT U5016 ( .A1(\read_value_mux[8][8] ), .A2(n1680), .A3(
        write_data[8]), .A4(n3092), .Y(\words[8]/data_i[8] ) );
  AO22X1_RVT U5017 ( .A1(\read_value_mux[8][9] ), .A2(n1680), .A3(
        write_data[9]), .A4(n3092), .Y(\words[8]/data_i[9] ) );
  AO21X1_RVT U5018 ( .A1(\words[8]/valid_o ), .A2(n1680), .A3(n3092), .Y(
        \words[8]/valid_i ) );
  AO22X1_RVT U5019 ( .A1(\read_value_mux[9][0] ), .A2(n1635), .A3(
        write_data[0]), .A4(n3097), .Y(\words[9]/data_i[0] ) );
  AO22X1_RVT U5020 ( .A1(\read_value_mux[9][10] ), .A2(n1635), .A3(
        write_data[10]), .A4(n3097), .Y(\words[9]/data_i[10] ) );
  AO22X1_RVT U5021 ( .A1(\read_value_mux[9][11] ), .A2(n1635), .A3(
        write_data[11]), .A4(n3097), .Y(\words[9]/data_i[11] ) );
  AO22X1_RVT U5022 ( .A1(\read_value_mux[9][12] ), .A2(n1635), .A3(
        write_data[12]), .A4(n3097), .Y(\words[9]/data_i[12] ) );
  AO22X1_RVT U5023 ( .A1(\read_value_mux[9][13] ), .A2(n1635), .A3(
        write_data[13]), .A4(n3097), .Y(\words[9]/data_i[13] ) );
  AO22X1_RVT U5024 ( .A1(\read_value_mux[9][14] ), .A2(n1635), .A3(
        write_data[14]), .A4(n3097), .Y(\words[9]/data_i[14] ) );
  AO22X1_RVT U5025 ( .A1(\read_value_mux[9][15] ), .A2(n1635), .A3(
        write_data[15]), .A4(n3097), .Y(\words[9]/data_i[15] ) );
  AO22X1_RVT U5026 ( .A1(\read_value_mux[9][16] ), .A2(n1635), .A3(
        write_data[16]), .A4(n3097), .Y(\words[9]/data_i[16] ) );
  AO22X1_RVT U5027 ( .A1(\read_value_mux[9][17] ), .A2(n1635), .A3(
        write_data[17]), .A4(n3097), .Y(\words[9]/data_i[17] ) );
  AO22X1_RVT U5028 ( .A1(\read_value_mux[9][18] ), .A2(n1635), .A3(
        write_data[18]), .A4(n3097), .Y(\words[9]/data_i[18] ) );
  AO22X1_RVT U5029 ( .A1(\read_value_mux[9][19] ), .A2(n1635), .A3(
        write_data[19]), .A4(n3097), .Y(\words[9]/data_i[19] ) );
  AO22X1_RVT U5030 ( .A1(\read_value_mux[9][1] ), .A2(n1635), .A3(
        write_data[1]), .A4(n3097), .Y(\words[9]/data_i[1] ) );
  AO22X1_RVT U5031 ( .A1(\read_value_mux[9][20] ), .A2(n1635), .A3(
        write_data[20]), .A4(n3097), .Y(\words[9]/data_i[20] ) );
  AO22X1_RVT U5032 ( .A1(\read_value_mux[9][21] ), .A2(n1635), .A3(
        write_data[21]), .A4(n3097), .Y(\words[9]/data_i[21] ) );
  AO22X1_RVT U5033 ( .A1(\read_value_mux[9][22] ), .A2(n1635), .A3(
        write_data[22]), .A4(n3097), .Y(\words[9]/data_i[22] ) );
  AO22X1_RVT U5034 ( .A1(\read_value_mux[9][23] ), .A2(n1635), .A3(
        write_data[23]), .A4(n3097), .Y(\words[9]/data_i[23] ) );
  AO22X1_RVT U5035 ( .A1(\read_value_mux[9][24] ), .A2(n1635), .A3(
        write_data[24]), .A4(n3097), .Y(\words[9]/data_i[24] ) );
  AO22X1_RVT U5036 ( .A1(\read_value_mux[9][25] ), .A2(n1635), .A3(
        write_data[25]), .A4(n3097), .Y(\words[9]/data_i[25] ) );
  AO22X1_RVT U5037 ( .A1(\read_value_mux[9][26] ), .A2(n1635), .A3(
        write_data[26]), .A4(n3097), .Y(\words[9]/data_i[26] ) );
  AO22X1_RVT U5038 ( .A1(\read_value_mux[9][27] ), .A2(n1635), .A3(
        write_data[27]), .A4(n3097), .Y(\words[9]/data_i[27] ) );
  AO22X1_RVT U5039 ( .A1(\read_value_mux[9][28] ), .A2(n1635), .A3(
        write_data[28]), .A4(n3097), .Y(\words[9]/data_i[28] ) );
  AO22X1_RVT U5040 ( .A1(\read_value_mux[9][29] ), .A2(n1635), .A3(
        write_data[29]), .A4(n3097), .Y(\words[9]/data_i[29] ) );
  AO22X1_RVT U5041 ( .A1(\read_value_mux[9][2] ), .A2(n1635), .A3(
        write_data[2]), .A4(n3097), .Y(\words[9]/data_i[2] ) );
  AO22X1_RVT U5042 ( .A1(n3097), .A2(write_data[30]), .A3(
        \read_value_mux[9][30] ), .A4(n1635), .Y(\words[9]/data_i[30] ) );
  AO22X1_RVT U5043 ( .A1(\read_value_mux[9][31] ), .A2(n1635), .A3(
        write_data[31]), .A4(n3097), .Y(\words[9]/data_i[31] ) );
  AO22X1_RVT U5044 ( .A1(\read_value_mux[9][3] ), .A2(n1635), .A3(
        write_data[3]), .A4(n3097), .Y(\words[9]/data_i[3] ) );
  AO22X1_RVT U5045 ( .A1(\read_value_mux[9][4] ), .A2(n1635), .A3(
        write_data[4]), .A4(n3097), .Y(\words[9]/data_i[4] ) );
  AO22X1_RVT U5046 ( .A1(\read_value_mux[9][5] ), .A2(n1635), .A3(
        write_data[5]), .A4(n3097), .Y(\words[9]/data_i[5] ) );
  AO22X1_RVT U5047 ( .A1(\read_value_mux[9][6] ), .A2(n1635), .A3(
        write_data[6]), .A4(n3097), .Y(\words[9]/data_i[6] ) );
  AO22X1_RVT U5048 ( .A1(\read_value_mux[9][7] ), .A2(n1635), .A3(
        write_data[7]), .A4(n3097), .Y(\words[9]/data_i[7] ) );
  AO22X1_RVT U5049 ( .A1(\read_value_mux[9][8] ), .A2(n1635), .A3(
        write_data[8]), .A4(n3097), .Y(\words[9]/data_i[8] ) );
  AO22X1_RVT U5050 ( .A1(\read_value_mux[9][9] ), .A2(n1635), .A3(
        write_data[9]), .A4(n3097), .Y(\words[9]/data_i[9] ) );
  AO21X1_RVT U5051 ( .A1(\words[9]/valid_o ), .A2(n1635), .A3(n3097), .Y(
        \words[9]/valid_i ) );
  NAND2X0_RVT U5052 ( .A1(n3112), .A2(n3111), .Y(n3113) );
endmodule

