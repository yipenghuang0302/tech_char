
module and_func ( a, b, y );
  input a, b;
  output y;


  AN2D0 U2 ( .A1(b), .A2(a), .Z(y) );
endmodule

